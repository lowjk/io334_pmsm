---------------------------------------------------------------------------------------------------------------------------------
-- Component name: PWM_OUTPUTPROTECTION
--
-- Synchronous: no 
--
-- Description: This component prevents A and B to be high at the exact same time. 
---------------------------------------------------------------------------------------------------------------------------------
 library IEEE; use IEEE.std_logic_1164.all; entity PWM_OUTPUTPROTECTION is port ( s0566B50C78A8B1778B34CE51EA1AE03DFB12AA1B : in std_logic_vector(1 downto 0); s6098D1E2037CC835C63EB95737225206F998214F : in std_logic; s529B64E065500EC35D88BFA7FDD85CEDD15C1CCD
 : in std_logic; s0D901D1A9772445D1277A56A33B3C8B7E4002BDF : out std_logic; s8A5BF12366BBF661A747D5AF98F670A7AC3B4888 : out std_logic ); end PWM_OUTPUTPROTECTION; architecture s44E7E05E235D0EE7F235C98FA35E8A7F01C7F087 of PWM_OUTPUTPROTECTION is constant s3E691753F846246E86D536A7B62303037FB148A4
 : std_logic_vector(1 downto 0) := "01"; constant sC87A65C9D0282A928184AA9652ABDFD6D576A746 : std_logic_vector(1 downto 0) := "10"; constant s44C5C6E4D8D98516A2EAFE9BCC864EA8911E21FF : std_logic_vector(1 downto 0) := "11"; begin      s0D901D1A9772445D1277A56A33B3C8B7E4002BDF
 <= '0' when s529B64E065500EC35D88BFA7FDD85CEDD15C1CCD = '1' and s0566B50C78A8B1778B34CE51EA1AE03DFB12AA1B = s3E691753F846246E86D536A7B62303037FB148A4 else '0' when s529B64E065500EC35D88BFA7FDD85CEDD15C1CCD = '1' and s0566B50C78A8B1778B34CE51EA1AE03DFB12AA1B
 = s44C5C6E4D8D98516A2EAFE9BCC864EA8911E21FF else s6098D1E2037CC835C63EB95737225206F998214F; s8A5BF12366BBF661A747D5AF98F670A7AC3B4888 <= '0' when s6098D1E2037CC835C63EB95737225206F998214F = '1' and s0566B50C78A8B1778B34CE51EA1AE03DFB12AA1B = sC87A65C9D0282A928184AA9652ABDFD6D576A746
 else '0' when s6098D1E2037CC835C63EB95737225206F998214F = '1' and s0566B50C78A8B1778B34CE51EA1AE03DFB12AA1B = s44C5C6E4D8D98516A2EAFE9BCC864EA8911E21FF else s529B64E065500EC35D88BFA7FDD85CEDD15C1CCD; end s44E7E05E235D0EE7F235C98FA35E8A7F01C7F087;