library IEEE; use IEEE.std_logic_1164.all; use IEEE.numeric_std.all; entity PWM_DELAY_ENABLE is port ( s82C78E3CD667612DE97ED7C5FA8365F21045093F : in std_logic; s0A61EC3B284D41A7527B973B71395AF396BD0749 : in std_logic; s90724AE20811A4A1CF4892AD6C5DE35913A379E1
 : in std_logic; s8198886663B13D3417529541102A2426672678BA : in std_logic_vector(31 downto 0); sE3594CA1813735566777C0F293E54987EE6AC901 : out std_logic ); end PWM_DELAY_ENABLE; architecture rtl of PWM_DELAY_ENABLE is signal s7BBA3C8AB08CE6CA89340ABD6C98D97CE084FAE3
, s12849FE6457414D598D01D43A97E8F0EB68AD8C6 : std_logic; signal s4EC95DE5C1C346B0D27A4875C7D0F0427B3047B4, s66943AE0205A978B8E4B0A809D118EF06B902F34 : unsigned(31 downto 0); begin process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749
) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749 = '1' then s4EC95DE5C1C346B0D27A4875C7D0F0427B3047B4 <= (others => '0'); elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then s4EC95DE5C1C346B0D27A4875C7D0F0427B3047B4 <= s66943AE0205A978B8E4B0A809D118EF06B902F34
; end if; end process; s66943AE0205A978B8E4B0A809D118EF06B902F34 <= s4EC95DE5C1C346B0D27A4875C7D0F0427B3047B4 + 1 when s90724AE20811A4A1CF4892AD6C5DE35913A379E1 = '1' else (others => '0'); process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749
) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749 = '1' then s7BBA3C8AB08CE6CA89340ABD6C98D97CE084FAE3 <= '0'; elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then s7BBA3C8AB08CE6CA89340ABD6C98D97CE084FAE3 <= s12849FE6457414D598D01D43A97E8F0EB68AD8C6
; end if; end process; s12849FE6457414D598D01D43A97E8F0EB68AD8C6 <= '0' when s90724AE20811A4A1CF4892AD6C5DE35913A379E1 = '0' else '1' when s90724AE20811A4A1CF4892AD6C5DE35913A379E1 = '1' and unsigned(s8198886663B13D3417529541102A2426672678BA) = 0 else '1' 
when s90724AE20811A4A1CF4892AD6C5DE35913A379E1 = '1' and s4EC95DE5C1C346B0D27A4875C7D0F0427B3047B4 = unsigned(s8198886663B13D3417529541102A2426672678BA) else s7BBA3C8AB08CE6CA89340ABD6C98D97CE084FAE3; sE3594CA1813735566777C0F293E54987EE6AC901 <= s7BBA3C8AB08CE6CA89340ABD6C98D97CE084FAE3
; end rtl;