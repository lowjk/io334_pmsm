library IEEE; use IEEE.std_logic_1164.all; entity PWM_EDGE_DETECTOR is port ( s82C78E3CD667612DE97ED7C5FA8365F21045093F : in std_logic; s0A61EC3B284D41A7527B973B71395AF396BD0749 : in std_logic; sAA3881E06E1AB1369AE662F6437029D7E01DC2A8 : in std_logic; s4EA41445886FECFF8F6DEA6BB5EB54DA56416129
 : out std_logic ); end PWM_EDGE_DETECTOR; architecture rtl of PWM_EDGE_DETECTOR is signal sDD1035FC1E341389045681CD6CD52DAA3469D282, sD9B608D5A96E68B773EBE94F8372AAE3B1EC7F52 : std_logic_vector(1 downto 0); begin process(s82C78E3CD667612DE97ED7C5FA8365F21045093F
, s0A61EC3B284D41A7527B973B71395AF396BD0749) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749 = '1' then sDD1035FC1E341389045681CD6CD52DAA3469D282 <= "00"; elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then sDD1035FC1E341389045681CD6CD52DAA3469D282
 <= sD9B608D5A96E68B773EBE94F8372AAE3B1EC7F52; end if; end process; sD9B608D5A96E68B773EBE94F8372AAE3B1EC7F52 <= sDD1035FC1E341389045681CD6CD52DAA3469D282(0) & sAA3881E06E1AB1369AE662F6437029D7E01DC2A8; s4EA41445886FECFF8F6DEA6BB5EB54DA56416129 <= '1' when
 sDD1035FC1E341389045681CD6CD52DAA3469D282 = "01" else '0'; end rtl;