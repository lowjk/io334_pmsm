library ieee; use ieee.std_logic_1164.all; package ENDAT_SNIFFER_pkg is  constant s731A256AA7EC109FE962BF102445534C5772925D : std_logic_vector(9 DOWNTO 0) := "00" & x"1B";  constant s7EC4167F3F7F1E99D074313BF18FF4BA05E7ED10 : std_logic_vector(9 DOWNTO 0) := "00" & x"01";
 constant s5907A17D8E29C7EB61D4F347241BFE4DAC407AEA : std_logic_vector(9 DOWNTO 0) := "00" & x"05";    constant sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81 : integer:= 6;  constant s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95 : integer:= 7;  constant s2B661762AEA08905D55D9C993A5A3B37FF2EC6CD
 : integer:= 32;  constant sCD3268FB2E69A058B357988C1BAD31C26B18C0D3 : integer:= 56;   constant sD086456116C26514BAA46126BDD5342689EA4666 : std_logic_vector(5 downto 0) := "000111";  constant sC950D600C869099649CD1A85609BA2714F805E57 : std_logic_vector(5 
downto 0) := "001110";  constant s37EC8A8DDC24DE5CCA325C6D520F09FE8B8BE3B0 : std_logic_vector(5 downto 0) := "011100";  constant sCE667A08F3FDC358AF7C3578CD6983F0DD93374C : std_logic_vector(5 downto 0) := "100011";  constant sEFA6395FD066E102662C9126CF88821C4940A5E2
 : std_logic_vector(5 downto 0) := "101010";  constant sA2C6EE455D0B31BBD6DC87409C4BCCEE5CFD35BD : std_logic_vector(5 downto 0) := "010101";  constant sBB116EDD54150FE461AF440792906CBAF166BCC9 : std_logic_vector(5 downto 0) := "110001";  constant s85EB2661C4F665AC828497B5A151BB556355E05B
 : std_logic_vector(5 downto 0) := "111000";  constant sAD320E17FE59D7A60E88C7BE1ADB0F57AA30EDD0 : std_logic_vector(5 downto 0) := "001001";  constant sA4D53F04E8BA4766E83AD0DEFDD9278B52C3044C : std_logic_vector(5 downto 0) := "011011";  constant sEDFBFD9F8F54F1BD9B20E33D40221B2D6C287A4D
 : std_logic_vector(5 downto 0) := "100100";  constant s9B0C1672B259D9C1E1031A2B01F0DF6FE98F2A2E : std_logic_vector(5 downto 0) := "101101";  constant sE78665F3E53F7F72C28BF19FCA20946AD4B10D08 : std_logic_vector(5 downto 0) := "110110";  constant s01C3860AF9A5F5F7A28F043ECA30EAB1DE4D786E
 : std_logic_vector(5 downto 0) := "010010";   function sC3DBD2E2D5E3454BB5656AA34F64BFD4C61C3377 (s6058A04FD298967655739A6C56676FA60DAE306B: in std_logic_vector) return std_logic_vector; end ENDAT_SNIFFER_pkg; package body ENDAT_SNIFFER_pkg is function sC3DBD2E2D5E3454BB5656AA34F64BFD4C61C3377
 (s6058A04FD298967655739A6C56676FA60DAE306B: in std_logic_vector) return std_logic_vector is variable s7CD850FFC99515521745FADBA902AC96D14969CA: std_logic_vector(s6058A04FD298967655739A6C56676FA60DAE306B'RANGE); alias sE8E6372BF4BD2203497CA7A3D999ACB746D3E75F
: std_logic_vector(s6058A04FD298967655739A6C56676FA60DAE306B'REVERSE_RANGE) is s6058A04FD298967655739A6C56676FA60DAE306B; begin for s020F5125771EEEB6F963720A8BB968FCA977AA41 in sE8E6372BF4BD2203497CA7A3D999ACB746D3E75F'RANGE loop s7CD850FFC99515521745FADBA902AC96D14969CA
(s020F5125771EEEB6F963720A8BB968FCA977AA41) := sE8E6372BF4BD2203497CA7A3D999ACB746D3E75F(s020F5125771EEEB6F963720A8BB968FCA977AA41); end loop; return s7CD850FFC99515521745FADBA902AC96D14969CA; end;  end ENDAT_SNIFFER_pkg; 