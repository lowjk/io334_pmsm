library ieee; use ieee.std_logic_1164.all; package ENDAT_ENCODER_memory_rom is  TYPE s3622567609DCA6521AA77BE1870D22909575B67D is array (integer range <>) of std_logic_vector(15 downto 0);  CONSTANT s1CFD18110A517486D9B5DAED3C58733F8D80465E : s3622567609DCA6521AA77BE1870D22909575B67D
(0 TO 1023) := (  X"0000",  X"0000",  X"0009",  X"10A9",   X"0000",  X"0000",  X"0000",  X"0000",  X"8003",  X"5053",  X"FF50",  X"FFFF",  X"50FF",  X"0000",  X"E001",  X"0000",   X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0001",  X"0000",  X"0000", 
 X"3031",  X"CD15",  X"075B",  X"B141",  X"DE68",  X"203A",  X"8000",  X"8001",   X"0800",  X"0401",  X"0104",  X"0000",  X"0000",  X"0029",  X"0000",  X"23E8",  X"3232",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"9873",   X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0E93",  X"4240",  X"000F",  X"0888",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",   X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0002", 
 X"3730",  X"3236",  X"3333",  X"0041",  X"6A63",  X"3277",  X"0000",  X"0001",  X"0000",  X"1420",  X"0000",  X"1420",  X"0000",  X"0001",  X"0000",  X"0001",  X"0000",  X"0001",  X"0000",  X"0001",  X"044C",  X"195A",  X"044C",  X"195A",  X"0000",  X"0001", 
 X"0258",  X"06EC",  X"0258",  X"06EC",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",   X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",   X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",   X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000"  );  CONSTANT sCD229F113F7E82913D1F47B1ED664487BEEB48A8 : s3622567609DCA6521AA77BE1870D22909575B67D(0 TO 1023) := (  X"000C",  X"0001", 
 X"0000",  X"8000",  X"8000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"FFFF",  X"FFFF",  X"FFFF",  X"FFFF",  X"0000",  X"8000",  X"494C",  X"3443",  X"3131",  X"2020",  X"0000",  X"0EF7",  X"0000",  X"0002",  X"1F40",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0800",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"8522",   X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",   X"000C",  X"0001",  X"0000",  X"8000",  X"8000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"FFFF",  X"FFFF",  X"FFFF",  X"FFFF",  X"0000",  X"8000",  X"494C",  X"3443",  X"3131",  X"2020",  X"0000",  X"0EF7",  X"0000",  X"0002",  X"1F40",  X"0000",  X"0000",  X"0000",  X"0000",  X"0800",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"8522",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000", 
 X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",  X"0000",   X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", 
 X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", 
 X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", 
 X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", 
 X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", 
 X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", 
 X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", 
 X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", 
 X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",  X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", 
 X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", 
 X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", 
 X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", 
 X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", 
 X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", 
 X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", 
 X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", 
 X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000" ); end ENDAT_ENCODER_memory_rom; 