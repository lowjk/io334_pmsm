library IEEE; use IEEE.std_logic_1164.all; use IEEE.numeric_std.all; entity PWM_DEADBAND is port ( s82C78E3CD667612DE97ED7C5FA8365F21045093F : in std_logic; s0A61EC3B284D41A7527B973B71395AF396BD0749 : in std_logic; sFE197AD05D9BDB6F66485EE431A46E7CAA1440DA
 : in std_logic_vector(15 downto 0); s4CEAF191FCC8603F876A2619B2DEE5520E94F8EB : in std_logic; sB3CC32098E3E0A09B7AE7118E531B3558C1C5529 : out std_logic ); end PWM_DEADBAND; architecture rtl of PWM_DEADBAND is type sA564510C7FCE7940D7D16C6D98FB4EC28EF9532B
 is (sCF4F5213523C5B43BD4A0FA51490511B11BDFB13, s778C688CC40AE12E8E4CA8998E4B784DE25AA00A); signal s0FEC712F765FB8844B3F2BBB11D39CEF1DC96CC4, s8E8B32351634161B9B1D8D18043D6DD1583B3BE6 : sA564510C7FCE7940D7D16C6D98FB4EC28EF9532B; signal s4F93C057303AA948FB806AB20CCA1F352C776944
, sB332F473DC201AE3FC8F7D31340A0D2F926BBE18 : std_logic_vector(1 downto 0); signal s669E87C26DAB148E4756B58CCB45860991766443 : std_logic; signal sE135D1BF1F08C5D8783FBC17D02365FB82575C41 : std_logic; signal sB22893CF06FAEE960448AD9991C03D88EB5846F7, s9EAF6EC1F95CED765E0651E3928D8B7CCB65372A
 : unsigned(15 downto 0); signal s011C53118C911BAD01FC70005A58267A477398BF : std_logic; signal s39D684145F6FD4C6D579F3BEC75102ECF4C39BAC : std_logic; signal s26FF4B7E9AE4046DC134099EAF5DB468745B34F9 : std_logic; begin    process(s82C78E3CD667612DE97ED7C5FA8365F21045093F
, s0A61EC3B284D41A7527B973B71395AF396BD0749) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749 = '1' then s4F93C057303AA948FB806AB20CCA1F352C776944 <= (others => '0'); elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then s4F93C057303AA948FB806AB20CCA1F352C776944
 <= sB332F473DC201AE3FC8F7D31340A0D2F926BBE18; end if; end process; sB332F473DC201AE3FC8F7D31340A0D2F926BBE18 <= s4F93C057303AA948FB806AB20CCA1F352C776944(0) & s4CEAF191FCC8603F876A2619B2DEE5520E94F8EB;  s669E87C26DAB148E4756B58CCB45860991766443 <= '1' when
 s4F93C057303AA948FB806AB20CCA1F352C776944 = "01" else '0';     process(s0FEC712F765FB8844B3F2BBB11D39CEF1DC96CC4, s669E87C26DAB148E4756B58CCB45860991766443, sFE197AD05D9BDB6F66485EE431A46E7CAA1440DA, sB22893CF06FAEE960448AD9991C03D88EB5846F7) begin  s011C53118C911BAD01FC70005A58267A477398BF
 <= '0'; s26FF4B7E9AE4046DC134099EAF5DB468745B34F9 <= '0'; s39D684145F6FD4C6D579F3BEC75102ECF4C39BAC <= '0'; case s0FEC712F765FB8844B3F2BBB11D39CEF1DC96CC4 is when sCF4F5213523C5B43BD4A0FA51490511B11BDFB13 => if s669E87C26DAB148E4756B58CCB45860991766443 = '1' 
then s011C53118C911BAD01FC70005A58267A477398BF <= '1'; s26FF4B7E9AE4046DC134099EAF5DB468745B34F9 <= '1'; s8E8B32351634161B9B1D8D18043D6DD1583B3BE6 <= s778C688CC40AE12E8E4CA8998E4B784DE25AA00A; else s8E8B32351634161B9B1D8D18043D6DD1583B3BE6 <= sCF4F5213523C5B43BD4A0FA51490511B11BDFB13
; end if; when s778C688CC40AE12E8E4CA8998E4B784DE25AA00A => if s669E87C26DAB148E4756B58CCB45860991766443 = '1' then s26FF4B7E9AE4046DC134099EAF5DB468745B34F9 <= '1'; s011C53118C911BAD01FC70005A58267A477398BF <= '1'; s8E8B32351634161B9B1D8D18043D6DD1583B3BE6
 <= s778C688CC40AE12E8E4CA8998E4B784DE25AA00A; elsif sB22893CF06FAEE960448AD9991C03D88EB5846F7 = unsigned(sFE197AD05D9BDB6F66485EE431A46E7CAA1440DA) then s26FF4B7E9AE4046DC134099EAF5DB468745B34F9 <= '1'; s011C53118C911BAD01FC70005A58267A477398BF <= '0'; s8E8B32351634161B9B1D8D18043D6DD1583B3BE6
 <= sCF4F5213523C5B43BD4A0FA51490511B11BDFB13; else s011C53118C911BAD01FC70005A58267A477398BF <= '1'; s39D684145F6FD4C6D579F3BEC75102ECF4C39BAC <= '1'; s8E8B32351634161B9B1D8D18043D6DD1583B3BE6 <= s778C688CC40AE12E8E4CA8998E4B784DE25AA00A; end if; end case
; end process; process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749 = '1' then s0FEC712F765FB8844B3F2BBB11D39CEF1DC96CC4 <= sCF4F5213523C5B43BD4A0FA51490511B11BDFB13
; elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then s0FEC712F765FB8844B3F2BBB11D39CEF1DC96CC4 <= s8E8B32351634161B9B1D8D18043D6DD1583B3BE6; end if; end process;     process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749
) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749 = '1' then sB22893CF06FAEE960448AD9991C03D88EB5846F7 <= (others => '0'); elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then sB22893CF06FAEE960448AD9991C03D88EB5846F7 <= s9EAF6EC1F95CED765E0651E3928D8B7CCB65372A
; end if; end process; s9EAF6EC1F95CED765E0651E3928D8B7CCB65372A <= (others => '0') when s26FF4B7E9AE4046DC134099EAF5DB468745B34F9 = '1' else sB22893CF06FAEE960448AD9991C03D88EB5846F7 + 1 when s39D684145F6FD4C6D579F3BEC75102ECF4C39BAC = '1' else sB22893CF06FAEE960448AD9991C03D88EB5846F7
;     sE135D1BF1F08C5D8783FBC17D02365FB82575C41 <= '0' when s011C53118C911BAD01FC70005A58267A477398BF = '1' else s4F93C057303AA948FB806AB20CCA1F352C776944(1);     sB3CC32098E3E0A09B7AE7118E531B3558C1C5529 <= s4F93C057303AA948FB806AB20CCA1F352C776944(1) when
 unsigned(sFE197AD05D9BDB6F66485EE431A46E7CAA1440DA) = 0 else sE135D1BF1F08C5D8783FBC17D02365FB82575C41; end rtl;