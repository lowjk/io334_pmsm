library IEEE; use IEEE.std_logic_1164.all; use IEEE.numeric_std.all; entity PWM_GENERATION is port ( s82C78E3CD667612DE97ED7C5FA8365F21045093F : in std_logic; s0A61EC3B284D41A7527B973B71395AF396BD0749 : in std_logic; s90724AE20811A4A1CF4892AD6C5DE35913A379E1
 : in std_logic; s67BC8086A3CA80A76AC4A164873CAD71C96B5FE0 : in std_logic_vector(7 downto 0); s160C88F52FE0264EE39CE02AD36940648A499C69 : in std_logic_vector(15 downto 0); s8AC4FA096044C5A37B22CAF70033FA5FE77D3BBA : in std_logic; s168C5AFF1BF7656559FC3937639C1AE2520B2927
 : in std_logic; s8FBFCA53F59AF345A2C3475B0AE37E3E7150F484 : in std_logic; sECA797D75838B39584026BAD00E0C439E8B77DD5 : in std_logic; sD246DF0225DF7A45E9F1ABE2CD12ADF9A529CE4F : in std_logic; s2C8B6CD97916AF6157800BCA22B0C2D46B5223EE : in std_logic; s37394BFF31F8165BDF20DEB888AECA974BBA3623
 : in std_logic_vector(31 downto 0); sBAF99F5E379DD83C7801574B6C9B3543793DAC97 : in std_logic_vector(31 downto 0); s210E8B1235B722AEADE3A804D3F0ABBF1ECDF813 : in std_logic_vector(31 downto 0); s3539C3439A2E15C9F92A30B0F8C66085F38548A7 : in std_logic_vector
(31 downto 0); s18DDC05E8E9DEDCDB9CE049E35C0239D9C743A48 : in std_logic_vector(31 downto 0); s503807568AF4A5E8CA829CD2CEE8004F3A340D32 : in std_logic_vector(31 downto 0); s933789B89707AE61A3E166FE17AA5F9396484D24 : in std_logic_vector(31 downto 0); s75E99097F31F71B794CA5D20959FA1D49963B501
 : out std_logic; s8A2ACBC26D8260C75D3D090B067684937C4AA807 : out std_logic; sB33828E1D3E6A13EBF56A658AFF3E791C2BCEF1D : out std_logic ); end PWM_GENERATION; architecture rtl of PWM_GENERATION is type sA564510C7FCE7940D7D16C6D98FB4EC28EF9532B is (sAD7CE844A8434A520DEEB9C7C1C7C0D7BCC9C3FA
, sBE4E204B6E36F17EA52DC2E02D321223132245AC); signal s0FEC712F765FB8844B3F2BBB11D39CEF1DC96CC4, s8E8B32351634161B9B1D8D18043D6DD1583B3BE6 : sA564510C7FCE7940D7D16C6D98FB4EC28EF9532B; signal s7EBC7B235873AE2953DA6A6511E8CB8F36CF4072, s21CECA1859128D26BA8CFD54FB491564917988EC
 : std_logic; signal s5DA1CF583D180062A64FE895478A6DC42F5C834C, sECED55B35F5E2505C16DDE8210E262A3CD4F2DAB : std_logic_vector(31 downto 0); signal s16D6ADEC9E8F6F1FDC56B50545E871AA893C9AC4, s7B22181EEF44DE728256FF0B191DBB5D3852E48A : std_logic_vector(31 downto
 0); signal sFE9F82A8AE8C792B89E09B771B1A919EE35E04EC, sCDA922F0F136064250C2A0B69C466CD0008B960F : std_logic_vector(31 downto 0); signal s99531FA05599F60BA2B3B189C8DD3E5C829863AD, s64A7755669160369452E1DF048419A8FAAD6A232 : unsigned(31 downto 0); signal sC336620F0A0095F6B6D6E13EAF03DA6990EAAC30
, s787C67DC96B4D37D71218A0C191895D5EF2EF824 : unsigned(31 downto 0); signal s4133DA6F31DC5E57FE03DEB9E8D54A257E8E629F, s7FC07F7407D6DD281CDD3D019FD095C3395DC863 : unsigned(31 downto 0); signal sBFFF49AD4F0F8DDD779E7A6AD18BAD7B76F69FD6 : std_logic_vector(31 
downto 0); signal s43D323C0CF5EABD478A64E350FC8F5B1DEE92488 : std_logic_vector(31 downto 0); signal s7FC0CF1421A8EDAC92B38A9018557B84F8F681E6 : std_logic; signal s323C9446EAAFB4A8E1D840DE84FE7BB7A1426FF4, s14DEA28292999031EA29E1B44A53236552DE0CE3 : unsigned
(31 downto 0); signal s9FE3AA951ED6F08B7A5413BDE7D4625290A5DE35, sFB21C382D397F043524483231D16DAD1BDAFFC78, sAF8B447761319CFA2D1422DE0ABB64BD107D5A00 : std_logic; signal s32EFBD3FB6C52E01480475AAAB3A00C2B0245F67 : std_logic; signal s66940A314138EA34FEDB71806200A98D45A20DAF
, s1DA93AF77962CDDA9A2F41296A6C97B1ED244E5C : std_logic; signal s74C20CCF9E09877336F0A793CC2883EEFEB474B9 : std_logic; signal s52CF23375D15A4333772E28BE7EAFDCD6C611361 : std_logic; signal s733A748A025F25F8E55BB915B70F4FE03871E777 : std_logic; signal sCA25B43014CB662A8D5E24A79A506675020AAFBC
 : std_logic; begin  sE801F5A846C27EDAD1E0D796BE9220AFD297BDF8: entity work.PWM_SHADOW port map ( s82C78E3CD667612DE97ED7C5FA8365F21045093F => s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749 => s0A61EC3B284D41A7527B973B71395AF396BD0749
, s5574F0669AE6133ED7FDB56FFBA9FE1BF90B7CA4 => s21CECA1859128D26BA8CFD54FB491564917988EC, s349EBE9125821C69A7A72BA275E6AFAF4C927A95 => s37394BFF31F8165BDF20DEB888AECA974BBA3623, sA5C3CFDDCDD135F575B15CDA6569B6A3284FA179 => s5DA1CF583D180062A64FE895478A6DC42F5C834C
 ); s82CAFED9C7D5F0F479614447710E71B7F7747BC9: entity work.PWM_SHADOW port map ( s82C78E3CD667612DE97ED7C5FA8365F21045093F => s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749 => s0A61EC3B284D41A7527B973B71395AF396BD0749
, s5574F0669AE6133ED7FDB56FFBA9FE1BF90B7CA4 => s21CECA1859128D26BA8CFD54FB491564917988EC, s349EBE9125821C69A7A72BA275E6AFAF4C927A95 => sBAF99F5E379DD83C7801574B6C9B3543793DAC97, sA5C3CFDDCDD135F575B15CDA6569B6A3284FA179 => sECED55B35F5E2505C16DDE8210E262A3CD4F2DAB
 ); s2C4A955E8A428E02DF441985E0BF5576BAA6490E: entity work.PWM_SHADOW port map ( s82C78E3CD667612DE97ED7C5FA8365F21045093F => s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749 => s0A61EC3B284D41A7527B973B71395AF396BD0749
, s5574F0669AE6133ED7FDB56FFBA9FE1BF90B7CA4 => s21CECA1859128D26BA8CFD54FB491564917988EC, s349EBE9125821C69A7A72BA275E6AFAF4C927A95 => s210E8B1235B722AEADE3A804D3F0ABBF1ECDF813, sA5C3CFDDCDD135F575B15CDA6569B6A3284FA179 => s16D6ADEC9E8F6F1FDC56B50545E871AA893C9AC4
 ); s47D83363D53E01C8A6A1AC48CB9119916E9B72B2: entity work.PWM_SHADOW port map ( s82C78E3CD667612DE97ED7C5FA8365F21045093F => s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749 => s0A61EC3B284D41A7527B973B71395AF396BD0749
, s5574F0669AE6133ED7FDB56FFBA9FE1BF90B7CA4 => s21CECA1859128D26BA8CFD54FB491564917988EC, s349EBE9125821C69A7A72BA275E6AFAF4C927A95 => s3539C3439A2E15C9F92A30B0F8C66085F38548A7, sA5C3CFDDCDD135F575B15CDA6569B6A3284FA179 => s7B22181EEF44DE728256FF0B191DBB5D3852E48A
 ); s67C2F61ADC856BFDC2AFBFAB8D26C2289FBD50F5: entity work.PWM_SHADOW port map ( s82C78E3CD667612DE97ED7C5FA8365F21045093F => s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749 => s0A61EC3B284D41A7527B973B71395AF396BD0749
, s5574F0669AE6133ED7FDB56FFBA9FE1BF90B7CA4 => s21CECA1859128D26BA8CFD54FB491564917988EC, s349EBE9125821C69A7A72BA275E6AFAF4C927A95 => s18DDC05E8E9DEDCDB9CE049E35C0239D9C743A48, sA5C3CFDDCDD135F575B15CDA6569B6A3284FA179 => sFE9F82A8AE8C792B89E09B771B1A919EE35E04EC
 ); sAEE68A85B77B1CFC3C4A56149761FB51F556EA74: entity work.PWM_SHADOW port map ( s82C78E3CD667612DE97ED7C5FA8365F21045093F => s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749 => s0A61EC3B284D41A7527B973B71395AF396BD0749
, s5574F0669AE6133ED7FDB56FFBA9FE1BF90B7CA4 => s21CECA1859128D26BA8CFD54FB491564917988EC, s349EBE9125821C69A7A72BA275E6AFAF4C927A95 => s503807568AF4A5E8CA829CD2CEE8004F3A340D32, sA5C3CFDDCDD135F575B15CDA6569B6A3284FA179 => sCDA922F0F136064250C2A0B69C466CD0008B960F
 ); s51F9E7A28AF8FA8E430A6B0E3C0D0B3C5B12ABEB: entity work.PWM_SHADOW port map ( s82C78E3CD667612DE97ED7C5FA8365F21045093F => s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749 => s0A61EC3B284D41A7527B973B71395AF396BD0749
, s5574F0669AE6133ED7FDB56FFBA9FE1BF90B7CA4 => s7EBC7B235873AE2953DA6A6511E8CB8F36CF4072,  s349EBE9125821C69A7A72BA275E6AFAF4C927A95 => s933789B89707AE61A3E166FE17AA5F9396484D24, sA5C3CFDDCDD135F575B15CDA6569B6A3284FA179 => sBFFF49AD4F0F8DDD779E7A6AD18BAD7B76F69FD6
 );  s43D323C0CF5EABD478A64E350FC8F5B1DEE92488 <= '0' & sBFFF49AD4F0F8DDD779E7A6AD18BAD7B76F69FD6(31 downto 1); s7FC0CF1421A8EDAC92B38A9018557B84F8F681E6 <= '1' when s323C9446EAAFB4A8E1D840DE84FE7BB7A1426FF4 = unsigned(s43D323C0CF5EABD478A64E350FC8F5B1DEE92488
) else '0'; s21CECA1859128D26BA8CFD54FB491564917988EC <= s7EBC7B235873AE2953DA6A6511E8CB8F36CF4072 or (s7FC0CF1421A8EDAC92B38A9018557B84F8F681E6 and sECA797D75838B39584026BAD00E0C439E8B77DD5) or sD246DF0225DF7A45E9F1ABE2CD12ADF9A529CE4F;      s9FE3AA951ED6F08B7A5413BDE7D4625290A5DE35
 <= '1' when unsigned(s5DA1CF583D180062A64FE895478A6DC42F5C834C) > unsigned(sECED55B35F5E2505C16DDE8210E262A3CD4F2DAB) else '0'; sFB21C382D397F043524483231D16DAD1BDAFFC78 <= '1' when unsigned(s16D6ADEC9E8F6F1FDC56B50545E871AA893C9AC4) > unsigned(s7B22181EEF44DE728256FF0B191DBB5D3852E48A
) else '0'; sAF8B447761319CFA2D1422DE0ABB64BD107D5A00 <= '1' when unsigned(sFE9F82A8AE8C792B89E09B771B1A919EE35E04EC) > unsigned(sCDA922F0F136064250C2A0B69C466CD0008B960F) else '0'; s99531FA05599F60BA2B3B189C8DD3E5C829863AD <= unsigned(s5DA1CF583D180062A64FE895478A6DC42F5C834C
) when s9FE3AA951ED6F08B7A5413BDE7D4625290A5DE35 = '0' else unsigned(sECED55B35F5E2505C16DDE8210E262A3CD4F2DAB); s64A7755669160369452E1DF048419A8FAAD6A232 <= unsigned(sECED55B35F5E2505C16DDE8210E262A3CD4F2DAB) when s9FE3AA951ED6F08B7A5413BDE7D4625290A5DE35
 = '0' else unsigned(s5DA1CF583D180062A64FE895478A6DC42F5C834C); sC336620F0A0095F6B6D6E13EAF03DA6990EAAC30 <= unsigned(s16D6ADEC9E8F6F1FDC56B50545E871AA893C9AC4) when sFB21C382D397F043524483231D16DAD1BDAFFC78 = '0' else unsigned(s7B22181EEF44DE728256FF0B191DBB5D3852E48A
); s787C67DC96B4D37D71218A0C191895D5EF2EF824 <= unsigned(s7B22181EEF44DE728256FF0B191DBB5D3852E48A) when sFB21C382D397F043524483231D16DAD1BDAFFC78 = '0' else unsigned(s16D6ADEC9E8F6F1FDC56B50545E871AA893C9AC4); s4133DA6F31DC5E57FE03DEB9E8D54A257E8E629F <= 
unsigned(sFE9F82A8AE8C792B89E09B771B1A919EE35E04EC) when sAF8B447761319CFA2D1422DE0ABB64BD107D5A00 = '0' else unsigned(sCDA922F0F136064250C2A0B69C466CD0008B960F); s7FC07F7407D6DD281CDD3D019FD095C3395DC863 <= unsigned(sCDA922F0F136064250C2A0B69C466CD0008B960F
) when sAF8B447761319CFA2D1422DE0ABB64BD107D5A00 = '0' else unsigned(sFE9F82A8AE8C792B89E09B771B1A919EE35E04EC);   process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749
 = '1' then s323C9446EAAFB4A8E1D840DE84FE7BB7A1426FF4 <= (others => '0'); elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then s323C9446EAAFB4A8E1D840DE84FE7BB7A1426FF4 <= s14DEA28292999031EA29E1B44A53236552DE0CE3; end if; end process; s14DEA28292999031EA29E1B44A53236552DE0CE3
 <= (others => '0') when s1DA93AF77962CDDA9A2F41296A6C97B1ED244E5C = '1' else s323C9446EAAFB4A8E1D840DE84FE7BB7A1426FF4 + 1 when s66940A314138EA34FEDB71806200A98D45A20DAF = '1' else s323C9446EAAFB4A8E1D840DE84FE7BB7A1426FF4; process(s0FEC712F765FB8844B3F2BBB11D39CEF1DC96CC4
, s323C9446EAAFB4A8E1D840DE84FE7BB7A1426FF4, sBFFF49AD4F0F8DDD779E7A6AD18BAD7B76F69FD6, s90724AE20811A4A1CF4892AD6C5DE35913A379E1, s2C8B6CD97916AF6157800BCA22B0C2D46B5223EE) begin  s32EFBD3FB6C52E01480475AAAB3A00C2B0245F67 <= '0'; s66940A314138EA34FEDB71806200A98D45A20DAF
 <= '0'; s1DA93AF77962CDDA9A2F41296A6C97B1ED244E5C <= '0'; s7EBC7B235873AE2953DA6A6511E8CB8F36CF4072 <= '0'; case s0FEC712F765FB8844B3F2BBB11D39CEF1DC96CC4 is when sAD7CE844A8434A520DEEB9C7C1C7C0D7BCC9C3FA => if s90724AE20811A4A1CF4892AD6C5DE35913A379E1 = '1' 
and s2C8B6CD97916AF6157800BCA22B0C2D46B5223EE = '0' then s1DA93AF77962CDDA9A2F41296A6C97B1ED244E5C <= '1'; s7EBC7B235873AE2953DA6A6511E8CB8F36CF4072 <= '1'; s8E8B32351634161B9B1D8D18043D6DD1583B3BE6 <= sBE4E204B6E36F17EA52DC2E02D321223132245AC; else s8E8B32351634161B9B1D8D18043D6DD1583B3BE6
 <= sAD7CE844A8434A520DEEB9C7C1C7C0D7BCC9C3FA; end if; when sBE4E204B6E36F17EA52DC2E02D321223132245AC => s32EFBD3FB6C52E01480475AAAB3A00C2B0245F67 <= '1'; if s323C9446EAAFB4A8E1D840DE84FE7BB7A1426FF4 = unsigned(sBFFF49AD4F0F8DDD779E7A6AD18BAD7B76F69FD6) then
 if s90724AE20811A4A1CF4892AD6C5DE35913A379E1 = '0' then s1DA93AF77962CDDA9A2F41296A6C97B1ED244E5C <= '1'; s8E8B32351634161B9B1D8D18043D6DD1583B3BE6 <= sAD7CE844A8434A520DEEB9C7C1C7C0D7BCC9C3FA; else s1DA93AF77962CDDA9A2F41296A6C97B1ED244E5C <= '1'; s7EBC7B235873AE2953DA6A6511E8CB8F36CF4072
 <= '1'; s8E8B32351634161B9B1D8D18043D6DD1583B3BE6 <= sBE4E204B6E36F17EA52DC2E02D321223132245AC; end if; elsif s2C8B6CD97916AF6157800BCA22B0C2D46B5223EE = '1' then s1DA93AF77962CDDA9A2F41296A6C97B1ED244E5C <= '1'; s8E8B32351634161B9B1D8D18043D6DD1583B3BE6
 <= sAD7CE844A8434A520DEEB9C7C1C7C0D7BCC9C3FA; else s66940A314138EA34FEDB71806200A98D45A20DAF <= '1'; s8E8B32351634161B9B1D8D18043D6DD1583B3BE6 <= sBE4E204B6E36F17EA52DC2E02D321223132245AC; end if; end case; end process; process(s82C78E3CD667612DE97ED7C5FA8365F21045093F
, s0A61EC3B284D41A7527B973B71395AF396BD0749) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749 = '1' then s0FEC712F765FB8844B3F2BBB11D39CEF1DC96CC4 <= sAD7CE844A8434A520DEEB9C7C1C7C0D7BCC9C3FA; elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) 
then s0FEC712F765FB8844B3F2BBB11D39CEF1DC96CC4 <= s8E8B32351634161B9B1D8D18043D6DD1583B3BE6; end if; end process;    s5B3C7C103E9F9155C1AD50978496F163C49FDA54: entity work.PWM_TRIGGER port map ( s82C78E3CD667612DE97ED7C5FA8365F21045093F => s82C78E3CD667612DE97ED7C5FA8365F21045093F
, s0A61EC3B284D41A7527B973B71395AF396BD0749 => s0A61EC3B284D41A7527B973B71395AF396BD0749, s4F9EF0C7BB9149A40FBFAFB249E3995FB864917A => s32EFBD3FB6C52E01480475AAAB3A00C2B0245F67, s67BC8086A3CA80A76AC4A164873CAD71C96B5FE0 => s67BC8086A3CA80A76AC4A164873CAD71C96B5FE0
, s96088CC8D215E1C4E6BD73028628BBAFD1FB4AB8 => std_logic_vector(s323C9446EAAFB4A8E1D840DE84FE7BB7A1426FF4), s160C88F52FE0264EE39CE02AD36940648A499C69 => s160C88F52FE0264EE39CE02AD36940648A499C69, s37394BFF31F8165BDF20DEB888AECA974BBA3623 => s5DA1CF583D180062A64FE895478A6DC42F5C834C
, sBAF99F5E379DD83C7801574B6C9B3543793DAC97 => sECED55B35F5E2505C16DDE8210E262A3CD4F2DAB, s210E8B1235B722AEADE3A804D3F0ABBF1ECDF813 => s16D6ADEC9E8F6F1FDC56B50545E871AA893C9AC4, s3539C3439A2E15C9F92A30B0F8C66085F38548A7 => s7B22181EEF44DE728256FF0B191DBB5D3852E48A
, s176765D58EB0F4B63A08449CD9D42334FA44A80B => (others => '0'), sFEE2B98E596E164B80FA91ED23A3B076B9EF6553 => s43D323C0CF5EABD478A64E350FC8F5B1DEE92488, sD570C51C1637403B1D115AC1158C653C42ECE9CB => s74C20CCF9E09877336F0A793CC2883EEFEB474B9 );    s52CF23375D15A4333772E28BE7EAFDCD6C611361
 <= '1' when (s323C9446EAAFB4A8E1D840DE84FE7BB7A1426FF4 >= s99531FA05599F60BA2B3B189C8DD3E5C829863AD) and (s323C9446EAAFB4A8E1D840DE84FE7BB7A1426FF4 < s64A7755669160369452E1DF048419A8FAAD6A232) and (s99531FA05599F60BA2B3B189C8DD3E5C829863AD /= s64A7755669160369452E1DF048419A8FAAD6A232
) else '0'; s733A748A025F25F8E55BB915B70F4FE03871E777 <= '1' when (s323C9446EAAFB4A8E1D840DE84FE7BB7A1426FF4 >= sC336620F0A0095F6B6D6E13EAF03DA6990EAAC30) and (s323C9446EAAFB4A8E1D840DE84FE7BB7A1426FF4 < s787C67DC96B4D37D71218A0C191895D5EF2EF824) and (sC336620F0A0095F6B6D6E13EAF03DA6990EAAC30
 /= s787C67DC96B4D37D71218A0C191895D5EF2EF824) else '0'; sCA25B43014CB662A8D5E24A79A506675020AAFBC <= '1' when (s323C9446EAAFB4A8E1D840DE84FE7BB7A1426FF4 >= s4133DA6F31DC5E57FE03DEB9E8D54A257E8E629F) and (s323C9446EAAFB4A8E1D840DE84FE7BB7A1426FF4 < s7FC07F7407D6DD281CDD3D019FD095C3395DC863
) and (s4133DA6F31DC5E57FE03DEB9E8D54A257E8E629F /= s7FC07F7407D6DD281CDD3D019FD095C3395DC863) else '0'; s75E99097F31F71B794CA5D20959FA1D49963B501 <= s8AC4FA096044C5A37B22CAF70033FA5FE77D3BBA when s32EFBD3FB6C52E01480475AAAB3A00C2B0245F67 = '0' else not s52CF23375D15A4333772E28BE7EAFDCD6C611361
 when s9FE3AA951ED6F08B7A5413BDE7D4625290A5DE35 = '1' else s52CF23375D15A4333772E28BE7EAFDCD6C611361; s8A2ACBC26D8260C75D3D090B067684937C4AA807 <= s168C5AFF1BF7656559FC3937639C1AE2520B2927 when s32EFBD3FB6C52E01480475AAAB3A00C2B0245F67 = '0' else not s733A748A025F25F8E55BB915B70F4FE03871E777
 when sFB21C382D397F043524483231D16DAD1BDAFFC78 = '1' else s733A748A025F25F8E55BB915B70F4FE03871E777; sB33828E1D3E6A13EBF56A658AFF3E791C2BCEF1D <= s8FBFCA53F59AF345A2C3475B0AE37E3E7150F484 when s32EFBD3FB6C52E01480475AAAB3A00C2B0245F67 = '0' else not (sCA25B43014CB662A8D5E24A79A506675020AAFBC
 or s74C20CCF9E09877336F0A793CC2883EEFEB474B9) when sAF8B447761319CFA2D1422DE0ABB64BD107D5A00 = '1' else sCA25B43014CB662A8D5E24A79A506675020AAFBC or s74C20CCF9E09877336F0A793CC2883EEFEB474B9; end rtl; 