library IEEE; use IEEE.STD_LOGIC_1164.all; entity PWM_SHADOW is PORT ( s82C78E3CD667612DE97ED7C5FA8365F21045093F : in std_logic; s0A61EC3B284D41A7527B973B71395AF396BD0749 : in std_logic; s5574F0669AE6133ED7FDB56FFBA9FE1BF90B7CA4 : in std_logic; s349EBE9125821C69A7A72BA275E6AFAF4C927A95
 : in std_logic_vector(31 downto 0); sA5C3CFDDCDD135F575B15CDA6569B6A3284FA179 : out std_logic_vector(31 downto 0) ); end PWM_SHADOW; architecture rtl of PWM_SHADOW is signal sF15ADA01195F0893D0DF096E72458BF060CAF275, sDF4D6BB37A0EADBB4FFF450A9A246DACDA52D258
 : std_logic_vector(31 downto 0); begin process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749 = '1' then sF15ADA01195F0893D0DF096E72458BF060CAF275 <= (others => '0'); elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then sF15ADA01195F0893D0DF096E72458BF060CAF275 <= sDF4D6BB37A0EADBB4FFF450A9A246DACDA52D258; end if; end process; sDF4D6BB37A0EADBB4FFF450A9A246DACDA52D258 <= s349EBE9125821C69A7A72BA275E6AFAF4C927A95
 when s5574F0669AE6133ED7FDB56FFBA9FE1BF90B7CA4 = '1' else sF15ADA01195F0893D0DF096E72458BF060CAF275; sA5C3CFDDCDD135F575B15CDA6569B6A3284FA179 <= sF15ADA01195F0893D0DF096E72458BF060CAF275; end rtl; 