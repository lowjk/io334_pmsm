--------------------------------------------------------------------------
-- Code Module version: 5
-- Why:
-- This PWM FPGA Code Module is intended to simplify much more the PWM
-- configuration.
-- PWM is high between On and Off.
--------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.PWM_pkg.all;

entity PWM is
  port
  (
    clk_i                      : in std_logic;
    reset_i                    : in std_logic;
    enable_i                   : in std_logic;
    idle_a_i                   : in std_logic;
    idle_b_i                   : in std_logic;
    idle_c_i                   : in std_logic;
    enable_latch_half_period_i : in std_logic;
    natural_pwm_update_i       : in std_logic;
    force_stop_i               : in std_logic;
    period_i                   : in std_logic_vector(31 downto 0);
    a_on_i                     : in std_logic_vector(31 downto 0);
    a_off_i                    : in std_logic_vector(31 downto 0);
    b_on_i                     : in std_logic_vector(31 downto 0);
    b_off_i                    : in std_logic_vector(31 downto 0);        
    c_on_i                     : in std_logic_vector(31 downto 0);
    c_off_i                    : in std_logic_vector(31 downto 0);
    deadband_i                 : in std_logic_vector(15 downto 0);
    protection_i               : in std_logic_vector( 1 downto 0);
    trigger_source_i           : in std_logic_vector( 7 downto 0);
    trigger_duration_i         : in std_logic_vector(15 downto 0);
    invert_a_i                 : in std_logic;
    invert_b_i                 : in std_logic;
    invert_c_i                 : in std_logic;
    version_o                  : out std_logic_vector(31 downto 0);
    delay_i                    : in std_logic_vector(31 downto 0);
    pwm_a_o                    : out std_logic;
    pwm_b_o                    : out std_logic;
    pwm_c_o                    : out std_logic
  );
end PWM;

  
architecture rtl of PWM is signal s52CF23375D15A4333772E28BE7EAFDCD6C611361, s733A748A025F25F8E55BB915B70F4FE03871E777, sCA25B43014CB662A8D5E24A79A506675020AAFBC : std_logic; signal sB1B3D4268C2B8B613C2FC8B041C841BAA0712B60, s6DB11F2CBC6D5D939FE7D2A0A15069F2CF271DA0
, s4FA28E14243B869FD010F952B61E89243E2BCBD5 : std_logic; signal s9188C71F17DB5E79F5E15D88BBC109099EA5C3D0, s13322D1A4BD74B670F14C8B0DC6A3541495F97B2 : std_logic; signal s7BBA3C8AB08CE6CA89340ABD6C98D97CE084FAE3 : std_logic; begin      s901AE81282F9EEA737FAA8F13EB1259D567DE2A6
: entity work.PWM_GENERATION port map ( s82C78E3CD667612DE97ED7C5FA8365F21045093F => clk_i, s0A61EC3B284D41A7527B973B71395AF396BD0749 => reset_i, s90724AE20811A4A1CF4892AD6C5DE35913A379E1 => s7BBA3C8AB08CE6CA89340ABD6C98D97CE084FAE3, s67BC8086A3CA80A76AC4A164873CAD71C96B5FE0
 => trigger_source_i, s160C88F52FE0264EE39CE02AD36940648A499C69 => trigger_duration_i, s8AC4FA096044C5A37B22CAF70033FA5FE77D3BBA => idle_a_i, s168C5AFF1BF7656559FC3937639C1AE2520B2927 => idle_b_i, s8FBFCA53F59AF345A2C3475B0AE37E3E7150F484 => idle_c_i, sECA797D75838B39584026BAD00E0C439E8B77DD5
 => enable_latch_half_period_i, sD246DF0225DF7A45E9F1ABE2CD12ADF9A529CE4F => natural_pwm_update_i, s2C8B6CD97916AF6157800BCA22B0C2D46B5223EE => force_stop_i, s37394BFF31F8165BDF20DEB888AECA974BBA3623 => a_on_i, sBAF99F5E379DD83C7801574B6C9B3543793DAC97 => 
a_off_i, s210E8B1235B722AEADE3A804D3F0ABBF1ECDF813 => b_on_i, s3539C3439A2E15C9F92A30B0F8C66085F38548A7 => b_off_i, s18DDC05E8E9DEDCDB9CE049E35C0239D9C743A48 => c_on_i, s503807568AF4A5E8CA829CD2CEE8004F3A340D32 => c_off_i, s933789B89707AE61A3E166FE17AA5F9396484D24
 => period_i, s75E99097F31F71B794CA5D20959FA1D49963B501 => s52CF23375D15A4333772E28BE7EAFDCD6C611361, s8A2ACBC26D8260C75D3D090B067684937C4AA807 => s733A748A025F25F8E55BB915B70F4FE03871E777, sB33828E1D3E6A13EBF56A658AFF3E791C2BCEF1D => sCA25B43014CB662A8D5E24A79A506675020AAFBC
 ); sF2EBA8E1D0F7D89614E1C708A4A8CCF27292D32A: entity work.PWM_DELAY_ENABLE port map ( s82C78E3CD667612DE97ED7C5FA8365F21045093F => clk_i, s0A61EC3B284D41A7527B973B71395AF396BD0749 => reset_i, s90724AE20811A4A1CF4892AD6C5DE35913A379E1 => enable_i, s8198886663B13D3417529541102A2426672678BA
 => delay_i, sE3594CA1813735566777C0F293E54987EE6AC901 => s7BBA3C8AB08CE6CA89340ABD6C98D97CE084FAE3 );           sC14ED7E869B04002F9FFB4995E3898FD1F9ED51D: entity work.PWM_DEADBAND port map ( s82C78E3CD667612DE97ED7C5FA8365F21045093F => clk_i, s0A61EC3B284D41A7527B973B71395AF396BD0749
 => reset_i, sFE197AD05D9BDB6F66485EE431A46E7CAA1440DA => deadband_i, s4CEAF191FCC8603F876A2619B2DEE5520E94F8EB => s52CF23375D15A4333772E28BE7EAFDCD6C611361, sB3CC32098E3E0A09B7AE7118E531B3558C1C5529 => sB1B3D4268C2B8B613C2FC8B041C841BAA0712B60 ); sFED8A944FE9E97B7F9282A1D168542B220E308FD
: entity work.PWM_DEADBAND port map ( s82C78E3CD667612DE97ED7C5FA8365F21045093F => clk_i, s0A61EC3B284D41A7527B973B71395AF396BD0749 => reset_i, sFE197AD05D9BDB6F66485EE431A46E7CAA1440DA => deadband_i, s4CEAF191FCC8603F876A2619B2DEE5520E94F8EB => s733A748A025F25F8E55BB915B70F4FE03871E777
, sB3CC32098E3E0A09B7AE7118E531B3558C1C5529 => s6DB11F2CBC6D5D939FE7D2A0A15069F2CF271DA0 );   s599AF2970DD5CE6F124431C571FA2FC04DC0F6DB: entity work.PWM_DEADBAND port map ( s82C78E3CD667612DE97ED7C5FA8365F21045093F => clk_i, s0A61EC3B284D41A7527B973B71395AF396BD0749
 => reset_i, sFE197AD05D9BDB6F66485EE431A46E7CAA1440DA => (others => '0'), s4CEAF191FCC8603F876A2619B2DEE5520E94F8EB => sCA25B43014CB662A8D5E24A79A506675020AAFBC, sB3CC32098E3E0A09B7AE7118E531B3558C1C5529 => s4FA28E14243B869FD010F952B61E89243E2BCBD5 );   
    sF734C4A48EE4DCBAF9ACD1CBC34E54EA143D9B2F: entity work.PWM_OUTPUTPROTECTION port map ( s0566B50C78A8B1778B34CE51EA1AE03DFB12AA1B => protection_i, s6098D1E2037CC835C63EB95737225206F998214F => sB1B3D4268C2B8B613C2FC8B041C841BAA0712B60, s529B64E065500EC35D88BFA7FDD85CEDD15C1CCD
 => s6DB11F2CBC6D5D939FE7D2A0A15069F2CF271DA0, s0D901D1A9772445D1277A56A33B3C8B7E4002BDF => s9188C71F17DB5E79F5E15D88BBC109099EA5C3D0, s8A5BF12366BBF661A747D5AF98F670A7AC3B4888 => s13322D1A4BD74B670F14C8B0DC6A3541495F97B2 );       version_o <= "10" & s731A256AA7EC109FE962BF102445534C5772925D
 & s7EC4167F3F7F1E99D074313BF18FF4BA05E7ED10 & s5907A17D8E29C7EB61D4F347241BFE4DAC407AEA; pwm_a_o <= not s9188C71F17DB5E79F5E15D88BBC109099EA5C3D0 when invert_a_i = '1' else s9188C71F17DB5E79F5E15D88BBC109099EA5C3D0; pwm_b_o <= not s13322D1A4BD74B670F14C8B0DC6A3541495F97B2
 when invert_b_i = '1' else s13322D1A4BD74B670F14C8B0DC6A3541495F97B2; pwm_c_o <= not s4FA28E14243B869FD010F952B61E89243E2BCBD5 when invert_c_i = '1' else s4FA28E14243B869FD010F952B61E89243E2BCBD5; end rtl; 