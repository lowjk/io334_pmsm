library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

  use work.BISS_ENCODER_pkg.all;

entity BISS_ENCODER is
  port
  (
    clk_i                 : in std_logic;
    reset_i               : in std_logic;
    
    version           : out std_logic_vector(31 downto 0); 
    
    busyDelay_i           : in std_logic_vector(31 downto 0); 
    lineDelay_i           : in std_logic_vector(9 downto 0);  
    numBits_i             : in std_logic_vector(7 downto 0);  
    timeoutClkCount_i     : in std_logic_vector(15 downto 0);      
    dataTxWord01_i        : in std_logic_vector(31 downto 0);
    dataTxWord02_i        : in std_logic_vector(31 downto 0);
    
    MA_i                  : in std_logic;
    SLI_i                 : in std_logic;  
    SLO_o                 : out std_logic
  );
end BISS_ENCODER;

architecture rtl of BISS_ENCODER is  signal s93E01125561FC324D133008782446ACFF4BEFAF7 : std_logic_vector(2 downto 0); signal sE61A76478B42ADEB9623894B73AED67882BFE166, s874E1C3DB6EE5D971219D07AF7042BDD48804660 : std_logic;  type sA564510C7FCE7940D7D16C6D98FB4EC28EF9532B
 is (s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C, sE0E4F2883171C2D3103F9C5E105BE2796C1D0D20, s4D0806694C40A4328E701B98C0CCFCF8D8018122, s0D68884FEE6B20EAD47E6890DB392A71177388C3, s04C04E81C51BCD79C38CAE4F767DB694E7C92F16, sB5ED9DCCE306B7A558C2A4CE5F0CE95BB735B7F1
, sB9C51836C6AC459392A2C47002628D79713F200E, s58B24B948EA83C487DAFFEC05D93C39626E147FF, s702D2C94BA354A47ED471B0C702D0BC853ED953A, sB26FAAB3194B59B57584637D1555B5E03B97A43E); signal sF1D6856D8C6E7F12EED89D6F5F90C7580EF3FE5E, sC3F360CDD6D534EE7E5EB80085F8A784CFE01687
 : sA564510C7FCE7940D7D16C6D98FB4EC28EF9532B;  signal sFB3107C8B48BCEDD631D98C6FE24FDE2FE5B35FC, s46222C520564F902D08A8F6AA78183FFD00C08A8 : std_logic; signal s1933CD31C2CAD7E35ECCFB532696A7E6679201C7 : unsigned(7 downto 0); signal s505B5BD52D1AB8AC55A87EE73A1FB0ADFEF658AD
, s8E67AEC73F44395450FB5D1F57AF753A7C92512E : std_logic; signal sCBF7EAA8073180E8522BAD491F6EF9A5E9803BFD : unsigned(31 downto 0); signal s785B9333AF11563F6096F3F423CD452D30979117 : std_logic; signal sA0F1804B53C834F4B3B21CBC401B64335F3ABD54 : std_logic; 
 signal s7D421768169CE02634C5F9A247D21A30EB3BA348 : unsigned(15 downto 0);  signal s5724103C905B1DD81E89674E48BBD9329E45720F : std_logic; signal sEA372DCD29AC0865067C5DA6367366307739297D : std_logic; signal s3011FB87583DAA89F74264003BDCBCD3B1AFD734 : std_logic_vector
(1023 downto 0); signal s0E8D465997071B21BE1B688F22BD23B325522377 : std_logic; signal s797CA649F8E0FFA9984E4E55CCD188314843F971 : std_logic_vector(63 downto 0); signal s3E30A5B3142B00CCBBD496C3953F892AFF63594A : integer range 0 to 63; begin version <= "10" & 
s731A256AA7EC109FE962BF102445534C5772925D & s7EC4167F3F7F1E99D074313BF18FF4BA05E7ED10 & s5907A17D8E29C7EB61D4F347241BFE4DAC407AEA;  s25EAD29E4C4980B19E612F54CC5B568B434EFE03: process(clk_i, reset_i) begin if reset_i = '1' then s93E01125561FC324D133008782446ACFF4BEFAF7
 <= (others => '0'); elsif rising_edge(clk_i) then s93E01125561FC324D133008782446ACFF4BEFAF7 <= s93E01125561FC324D133008782446ACFF4BEFAF7(1 downto 0) & MA_i; end if; end process s25EAD29E4C4980B19E612F54CC5B568B434EFE03; sE61A76478B42ADEB9623894B73AED67882BFE166
 <= '1' when s93E01125561FC324D133008782446ACFF4BEFAF7(2 downto 1) = "01" else '0'; s874E1C3DB6EE5D971219D07AF7042BDD48804660 <= '1' when s93E01125561FC324D133008782446ACFF4BEFAF7(2 downto 1) = "10" else '0';  sA0E3F628288F9FF5ED44D93BDADE0807C5D95734 : process
(sF1D6856D8C6E7F12EED89D6F5F90C7580EF3FE5E, s874E1C3DB6EE5D971219D07AF7042BDD48804660, sE61A76478B42ADEB9623894B73AED67882BFE166, sCBF7EAA8073180E8522BAD491F6EF9A5E9803BFD, busyDelay_i, s1933CD31C2CAD7E35ECCFB532696A7E6679201C7, numBits_i, s7D421768169CE02634C5F9A247D21A30EB3BA348
, timeoutClkCount_i, sEA372DCD29AC0865067C5DA6367366307739297D, s785B9333AF11563F6096F3F423CD452D30979117) begin  s0E8D465997071B21BE1B688F22BD23B325522377 <= '1'; s505B5BD52D1AB8AC55A87EE73A1FB0ADFEF658AD <= '0'; sFB3107C8B48BCEDD631D98C6FE24FDE2FE5B35FC
 <= '0'; s8E67AEC73F44395450FB5D1F57AF753A7C92512E <= '0'; s46222C520564F902D08A8F6AA78183FFD00C08A8 <= '0'; s5724103C905B1DD81E89674E48BBD9329E45720F <= '0'; sA0F1804B53C834F4B3B21CBC401B64335F3ABD54 <= '0'; case sF1D6856D8C6E7F12EED89D6F5F90C7580EF3FE5E
 is when s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C => s0E8D465997071B21BE1B688F22BD23B325522377 <= '1'; s505B5BD52D1AB8AC55A87EE73A1FB0ADFEF658AD <= '1'; sFB3107C8B48BCEDD631D98C6FE24FDE2FE5B35FC <= '1'; sA0F1804B53C834F4B3B21CBC401B64335F3ABD54 <= '1'; if
 s874E1C3DB6EE5D971219D07AF7042BDD48804660 ='1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= sE0E4F2883171C2D3103F9C5E105BE2796C1D0D20; else sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C; end if; when sE0E4F2883171C2D3103F9C5E105BE2796C1D0D20
 => s0E8D465997071B21BE1B688F22BD23B325522377 <= '1'; s5724103C905B1DD81E89674E48BBD9329E45720F <= '1'; if sE61A76478B42ADEB9623894B73AED67882BFE166 = '1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s4D0806694C40A4328E701B98C0CCFCF8D8018122; elsif s785B9333AF11563F6096F3F423CD452D30979117
 = '1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C; else sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= sE0E4F2883171C2D3103F9C5E105BE2796C1D0D20; end if; when s4D0806694C40A4328E701B98C0CCFCF8D8018122 => s0E8D465997071B21BE1B688F22BD23B325522377
 <= '1'; if sE61A76478B42ADEB9623894B73AED67882BFE166 = '1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s0D68884FEE6B20EAD47E6890DB392A71177388C3; elsif s785B9333AF11563F6096F3F423CD452D30979117 = '1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= 
s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C; else sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s4D0806694C40A4328E701B98C0CCFCF8D8018122; end if; when s0D68884FEE6B20EAD47E6890DB392A71177388C3 => s0E8D465997071B21BE1B688F22BD23B325522377 <= '0'; s8E67AEC73F44395450FB5D1F57AF753A7C92512E
 <= '1'; if sCBF7EAA8073180E8522BAD491F6EF9A5E9803BFD >= unsigned(busyDelay_i) then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s04C04E81C51BCD79C38CAE4F767DB694E7C92F16; else sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s0D68884FEE6B20EAD47E6890DB392A71177388C3
; end if; when s04C04E81C51BCD79C38CAE4F767DB694E7C92F16 => s0E8D465997071B21BE1B688F22BD23B325522377 <= '0'; if sE61A76478B42ADEB9623894B73AED67882BFE166 = '1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= sB5ED9DCCE306B7A558C2A4CE5F0CE95BB735B7F1; elsif
 s785B9333AF11563F6096F3F423CD452D30979117 = '1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C; else sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s04C04E81C51BCD79C38CAE4F767DB694E7C92F16; end if; when sB5ED9DCCE306B7A558C2A4CE5F0CE95BB735B7F1
 => s0E8D465997071B21BE1B688F22BD23B325522377 <= '1'; if sE61A76478B42ADEB9623894B73AED67882BFE166 = '1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= sB9C51836C6AC459392A2C47002628D79713F200E; elsif s785B9333AF11563F6096F3F423CD452D30979117 = '1' then
 sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C; else sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= sB5ED9DCCE306B7A558C2A4CE5F0CE95BB735B7F1; end if; when sB9C51836C6AC459392A2C47002628D79713F200E => s0E8D465997071B21BE1B688F22BD23B325522377
 <= '0'; if sE61A76478B42ADEB9623894B73AED67882BFE166 = '1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s58B24B948EA83C487DAFFEC05D93C39626E147FF; elsif s785B9333AF11563F6096F3F423CD452D30979117 = '1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= 
s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C; else sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= sB9C51836C6AC459392A2C47002628D79713F200E; end if; when s58B24B948EA83C487DAFFEC05D93C39626E147FF => s0E8D465997071B21BE1B688F22BD23B325522377 <= sEA372DCD29AC0865067C5DA6367366307739297D
; if sE61A76478B42ADEB9623894B73AED67882BFE166 = '1' and s1933CD31C2CAD7E35ECCFB532696A7E6679201C7 < unsigned(numBits_i)-1 then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s702D2C94BA354A47ED471B0C702D0BC853ED953A; elsif sE61A76478B42ADEB9623894B73AED67882BFE166
 = '1' and s1933CD31C2CAD7E35ECCFB532696A7E6679201C7 >= unsigned(numBits_i)-1 then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= sB26FAAB3194B59B57584637D1555B5E03B97A43E; elsif s785B9333AF11563F6096F3F423CD452D30979117 = '1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687
 <= s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C; else sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s58B24B948EA83C487DAFFEC05D93C39626E147FF; end if; when s702D2C94BA354A47ED471B0C702D0BC853ED953A => s0E8D465997071B21BE1B688F22BD23B325522377 <= sEA372DCD29AC0865067C5DA6367366307739297D
; s46222C520564F902D08A8F6AA78183FFD00C08A8 <= '1'; sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s58B24B948EA83C487DAFFEC05D93C39626E147FF; when sB26FAAB3194B59B57584637D1555B5E03B97A43E => s0E8D465997071B21BE1B688F22BD23B325522377 <= '0'; if s785B9333AF11563F6096F3F423CD452D30979117
 = '1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C; else sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= sB26FAAB3194B59B57584637D1555B5E03B97A43E; end if; end case; end process sA0E3F628288F9FF5ED44D93BDADE0807C5D95734
;  s01B836CC599AAC170C41C635FD46B72FA2B88119: process(clk_i, reset_i) begin if reset_i = '1' then sF1D6856D8C6E7F12EED89D6F5F90C7580EF3FE5E <= s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C; elsif rising_edge(clk_i) then sF1D6856D8C6E7F12EED89D6F5F90C7580EF3FE5E
 <= sC3F360CDD6D534EE7E5EB80085F8A784CFE01687; end if; end process s01B836CC599AAC170C41C635FD46B72FA2B88119;  s3B22EB14E3B344A665CDCFA537682F683F817270: process(clk_i, reset_i) begin if reset_i = '1' then sCBF7EAA8073180E8522BAD491F6EF9A5E9803BFD <= (others
 => '0'); elsif rising_edge(clk_i) then if s505B5BD52D1AB8AC55A87EE73A1FB0ADFEF658AD = '1' then sCBF7EAA8073180E8522BAD491F6EF9A5E9803BFD <= (others => '0'); elsif s8E67AEC73F44395450FB5D1F57AF753A7C92512E='1' then sCBF7EAA8073180E8522BAD491F6EF9A5E9803BFD
 <= sCBF7EAA8073180E8522BAD491F6EF9A5E9803BFD + 1; end if; end if; end process s3B22EB14E3B344A665CDCFA537682F683F817270;  sE89B484851192CC4812859B8C19EB7C1BC90F325: process(clk_i, reset_i) begin if reset_i = '1' then s7D421768169CE02634C5F9A247D21A30EB3BA348
 <= (others => '0'); s785B9333AF11563F6096F3F423CD452D30979117 <= '0'; elsif rising_edge(clk_i) then if sE61A76478B42ADEB9623894B73AED67882BFE166='1' or s874E1C3DB6EE5D971219D07AF7042BDD48804660='1' then s7D421768169CE02634C5F9A247D21A30EB3BA348 <= (others
 => '0'); s785B9333AF11563F6096F3F423CD452D30979117 <= '0'; elsif s7D421768169CE02634C5F9A247D21A30EB3BA348 < unsigned(timeOutClkCount_i) then s7D421768169CE02634C5F9A247D21A30EB3BA348 <= s7D421768169CE02634C5F9A247D21A30EB3BA348 + 1; s785B9333AF11563F6096F3F423CD452D30979117
 <= '0'; else s785B9333AF11563F6096F3F423CD452D30979117 <= '1'; end if; end if; end process sE89B484851192CC4812859B8C19EB7C1BC90F325;  sE96D7A9A7A11F700AE10FCF23B2615B196036470: process(clk_i, reset_i) begin if reset_i = '1' then s3011FB87583DAA89F74264003BDCBCD3B1AFD734
 <= (others => '1'); elsif rising_edge(clk_i) then if sA0F1804B53C834F4B3B21CBC401B64335F3ABD54='1' then s3011FB87583DAA89F74264003BDCBCD3B1AFD734 <= (others => '1'); else s3011FB87583DAA89F74264003BDCBCD3B1AFD734 <= s3011FB87583DAA89F74264003BDCBCD3B1AFD734
(1022 downto 0) & s0E8D465997071B21BE1B688F22BD23B325522377; end if; end if; end process sE96D7A9A7A11F700AE10FCF23B2615B196036470; s04F1C1995ECB20E1F71B35E2D1D3AFA2C11F71CC : process(lineDelay_i, s3011FB87583DAA89F74264003BDCBCD3B1AFD734) begin for s020F5125771EEEB6F963720A8BB968FCA977AA41
 in 0 to 1023 loop if s020F5125771EEEB6F963720A8BB968FCA977AA41=to_integer(unsigned(lineDelay_i)) then SLO_o <= s3011FB87583DAA89F74264003BDCBCD3B1AFD734(s020F5125771EEEB6F963720A8BB968FCA977AA41); end if; end loop; end process s04F1C1995ECB20E1F71B35E2D1D3AFA2C11F71CC
;  s1A6B9D64C1C1642B9CE9DAD04D5D0F4EE65A3846: process(clk_i, reset_i) begin if reset_i = '1' then s797CA649F8E0FFA9984E4E55CCD188314843F971 <= (others => '0'); elsif rising_edge(clk_i) then if s5724103C905B1DD81E89674E48BBD9329E45720F = '1' then s797CA649F8E0FFA9984E4E55CCD188314843F971
 <= dataTxWord02_i & dataTxWord01_i; end if; end if; end process s1A6B9D64C1C1642B9CE9DAD04D5D0F4EE65A3846;  s3E30A5B3142B00CCBBD496C3953F892AFF63594A <= to_integer(unsigned(numBits_i)-s1933CD31C2CAD7E35ECCFB532696A7E6679201C7-1); sEC722CF0BB8881E6BBF8D954FCA31E95819A3196
 : process(numBits_i, s1933CD31C2CAD7E35ECCFB532696A7E6679201C7, s797CA649F8E0FFA9984E4E55CCD188314843F971, s3E30A5B3142B00CCBBD496C3953F892AFF63594A) begin for s020F5125771EEEB6F963720A8BB968FCA977AA41 in 0 to 63 loop if s020F5125771EEEB6F963720A8BB968FCA977AA41
=s3E30A5B3142B00CCBBD496C3953F892AFF63594A then sEA372DCD29AC0865067C5DA6367366307739297D <= s797CA649F8E0FFA9984E4E55CCD188314843F971(s020F5125771EEEB6F963720A8BB968FCA977AA41); end if; end loop; end process sEC722CF0BB8881E6BBF8D954FCA31E95819A3196;  s28878808207CD2A29EA2B709A742EB4D419FA7CF
: process(clk_i, reset_i) begin if reset_i = '1' then s1933CD31C2CAD7E35ECCFB532696A7E6679201C7 <= (others => '0'); elsif rising_edge(clk_i) then if sFB3107C8B48BCEDD631D98C6FE24FDE2FE5B35FC = '1' then s1933CD31C2CAD7E35ECCFB532696A7E6679201C7 <= (others => '0'); elsif s46222C520564F902D08A8F6AA78183FFD00C08A8 = '1' then s1933CD31C2CAD7E35ECCFB532696A7E6679201C7 <= s1933CD31C2CAD7E35ECCFB532696A7E6679201C7 + 1; end if; end if; end process s28878808207CD2A29EA2B709A742EB4D419FA7CF; end rtl;