library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;
  use work.ENDAT_ENCODER_pkg.all;
  use work.ENDAT_ENCODER_memory_rom.all;

entity ENDAT_ENCODER is
  port
  (
    clk_i            : in std_logic;
    reset_i          : in std_logic;

    
    version_o        : out std_logic_vector(31 downto 0);

    
    td_i             : in std_logic_vector(31 downto 0);  
    tm_i             : in std_logic_vector(31 downto 0);  
    tR_i             : in std_logic_vector(31 downto 0);  
    tcal_i           : in std_logic_vector(31 downto 0);  
    numPulPosVal_i   : in std_logic_vector(31 downto 0);  
    distRev_i        : in std_logic_vector(31 downto 0);  
    temperature_i    : in std_logic_vector(31 downto 0);
    commutation_i    : in std_logic_vector(31 downto 0);

    
    dataMode_i       : in std_logic_vector(31 downto 0);  
    dataRx_LSB_i     : in std_logic_vector(31 downto 0);  
    dataRx_MSB_i     : in std_logic_vector(31 downto 0);  

    
    o_serial      : out std_logic;  
    i_serial_clk  : in std_logic;   
    i_serial      : in std_logic;   
    o_drive_en    : out std_logic   
  );
end ENDAT_ENCODER;

architecture Struct OF ENDAT_ENCODER IS   constant sED14BC4B3908B6DB77B3D546FFC4257CF3675A4F : std_logic := '1'; constant sC74718EA1B32E1BE7F9362F1CB8194555A8B7321 : unsigned(31 downto 0) := to_unsigned( 2, 32); constant sC1671CA18999DFAA45150AF19CC9FCDC05B45FC2
 : unsigned(31 downto 0) := to_unsigned( 6, 32); constant s73B96A69A181F16E9161FFCBBB71691BE5986214 : unsigned(31 downto 0) := to_unsigned( 8, 32); constant s0C8BF396CD56CBB5C916487998FFF3E0646F0DA8 : unsigned(31 downto 0) := to_unsigned(16, 32); constant
 sAC85A76D3768A4693698919CFE1AC38E3EC7E60B : unsigned(31 downto 0) := to_unsigned( 3, 32); constant s7F754F692527BC0267C69BBEFF22B0EB623D725D : unsigned(31 downto 0) := to_unsigned( 8, 32); constant sE417F33BECFBA77833DA36525F430E5AEB7C96D5 : unsigned(31 
downto 0) := to_unsigned(30, 32);   constant sD0F92C1D45611463356A15CFF87B99280A8A24F1 : unsigned(21 downto 0) := to_unsigned( 594000,22);  constant sB6C4B6996BE4000D3F7E6A44BB9ED1B6A592CAF0 : unsigned(21 downto 0) := to_unsigned( 65536,22);  constant s2E3247119760310EEBE0E32A775CFE4D34F8DD21
 : unsigned( 3 downto 0) := to_unsigned( 8, 4);  constant s180C3B3A658D0B94ADDD3EBA8B3FD02288454264 : unsigned( 3 downto 0) := to_unsigned( 10, 4);  constant s768F8BF346D525F17E3ACF7560EB0D135C6F4041 : unsigned(21 downto 0) := to_unsigned(3750938,22);    
 type sCBF5A8DB3DE001E3C6479CF4BC6B0BE6407CA993 is (s4EEF46B8032D06418C2A950FC6E48D5A56D77264, sBB12D33790A5D3018B4D986F4ADB83977C5D8601, s39392447A31070974A90414173657878F7BACB37, s80DC381C4925691B4334DD614AE199EF1D448C52, s67E7CF8001D8C888E6037A63B2A88D9E50C20BF3
, sED64C84C9A97C77A28959EB3D8FD87CFD05499E0, sC8D8E0168DF0925533D8199135EDFCE49E855CE9, s58B24B948EA83C487DAFFEC05D93C39626E147FF, s88BB3E464A5433B5E70C481850CFB4250671F723, s13CF374CF3BFFB5D28DC3FA96C2EDB6E5F3847E9, sB75F5ECEEDFEADF68941469BEA18B3230DC55E12
, sC9891EDB20266FE6D4FB2432877D93C6F27E651B, s9361618BB4D0D11E48353A207CDF79F17E90ECC6, sD1A28D5936291214869D8F06C0ADAF373A1B02C6, s1375AEE1631E1F16F7F548230C9A174D991B8343, s51B97BD443CF4AC466F639B508697B38106C2BA3, s46DB2160F9823D6161D8CD94822C414FA337C670
, sE39C1BB78C737B4D4A9AEC7FAE586981C1DD6B52);  type s742C0B6CE6500669B746A3B43B9F603B1E3EE0D3 is (s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C, s89180489BEBF665610DC5098AB8F99C0BBF612FE, sF0D99209603F6F7473DE58A048ABB74800BF9B6E, sB72BA5545AAD812117645A3F42558C3927D9E971
, sE73FCB3053E16A73428686A101357781139D2C9D, s0FC3DA9494BAFC3ED1F299DDF23029966E219F55);    signal s39BBA73E802D1EC6F9481E64A0C553405F91F14A : std_logic_vector(1 to 3) := (others => '0'); signal s1BACD241F56E4F52722832FA830845B2068BC767, s03C86E6A8EC0C1604AE1C69CEB6A81B140CF163E
 : std_logic; signal sDD66F717A56E6D482292350AFE88447E9E2FB37F : std_logic_vector(1 to 2) := (others => '0'); signal s5C9DDF5B777BD5A3F655299884019D187CEB0736 : std_logic := '0'; signal s5195EFEEEF3FA327D997E7C77C21627F37E4F83C : std_logic;  signal s7437C738E80B44EBF7CA42B918E6968B6656249F
, s5FDA25AB9BF862813FA68F7621B5928C66206883 : sCBF5A8DB3DE001E3C6479CF4BC6B0BE6407CA993;  signal s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E : std_logic_vector( 5 downto 0) := (others => '0'); signal sD379CAE4835BBA8234DDEC3E02227FC8A456159E : std_logic_vector
( 7 downto 0) := (others => '0'); signal sCDC84BF1C2EA12755C5188D514BC2D52B0FD0981 : std_logic_vector(15 downto 0) := (others => '0');  signal s74479D486ED1C3DA5D4D8F982E552DE6F4019633 : std_logic_vector(7 downto 0) := (others => '0'); signal s49778255829DFE971575864AE71D03CF1A0C4867
 : std_logic_vector(7 downto 0) := (others => '0'); signal s10C1DD445A18FDB20BE62ADD7A9A8635E879AD33 : std_logic_vector(7 downto 0) := s57E60BF34E25CCC564142C57DBFF63876615DB5E; signal sF74B9451531F47DEF952886360EE46EDA03FABA6 : std_logic_vector(7 downto 0) := 
s83F243E9AEA0950EEEE87EEFF9FF2B8AA0412294;  signal s1E02444D182262D00D4A327664194E0E7C9BCD58, s61E8DE0133C8A0EA7C46D3E5F1005799218FEF8B : s742C0B6CE6500669B746A3B43B9F603B1E3EE0D3; signal s440318DC9344B28FB76FFB67D03C27AF3B02548D : std_logic; signal sF4A7A88B0CE794196EC3287991182494C4CF68BB
 : std_logic;  signal sFF8DA13899BDB1FC1B166E7DBE024EA19D9D8E78 : unsigned( 3 downto 0) := (others => '0'); signal sFD38B58449B1F8FD27CEFABE026072920D7C6664 : unsigned(21 downto 0) := (others => '0'); signal s3E66115776824191EC46FFEDCE8964F683B11326 : unsigned
( 5 downto 0) := (others => '0'); signal sBCFB815ECFC1ADE1DD3A8C00366D0325652CDF68 : unsigned(21 downto 0) := (others => '0'); signal s34682EDE73B453730FDDB73AE693BF6858792888 : unsigned(15 downto 0) := (others => '0'); signal s8A2992E6D362DBB70C96CD6B71F48399524E30D2
 : unsigned(21 downto 0) := (others => '0');  signal s0399AD38FFE6E9911310CCF2C7975E26207D5D3D : integer range 0 to 63; signal sAABA4D54E9D1D3E0E35625A7E9DAF3FECB7C633F : unsigned(5 downto 0); signal sD2575E546E2EC143C5C4DD4FCD988505DC92A552 : std_logic_vector
(47 downto 0); signal sCFD226CC0ECDD9D07EE7E693ABB8A3A3B1E2CF73 : std_logic_vector(47 downto 0); signal sEE8C5684D6E32E443D201C83D1FDFBBBAC150FAD : std_logic_vector(47 downto 0); signal sC4B6EA407C3AA8DD2E6A18E7F77C14FACC951414, s06E676C0BDF7C68FD7495790A14A2FEBA13D3DB6
, warning, s76804DD01BB29A387010BCE68256FDB2A4020735, sCB42C2FDABBD75F13A77BB4E139059E0A23744FD : std_logic; signal sBB999F79F35F7555095A7373986DE0689DE5FC46 : std_logic_vector(50 downto 0); signal sEF80C7392E78A56484621A1127C5B6AB5F281091 : std_logic_vector
(24 downto 0); signal sDDFA38A34F7901FE6E261DE887A8F537753CF545 : std_logic_vector(24 downto 0);  signal sAE11F5A23788CBD8FAF306A52CAC70458125557A : std_logic_vector(50 downto 0) := (others => '0'); signal sCFF2D518C744D824B9DE2B4D9AFBF5F4725457B2 : std_logic_vector
(24 downto 0) := (others => '0'); signal sB355DE414F49CCFFF6381B960907D94AA7FBF024 : std_logic_vector(24 downto 0) := (others => '0'); signal s63B7F7C57F075889730F3ADD94597ABD229977FB : std_logic_vector(4 downto 0) := (others => '1'); signal sD3C21919EB55E97996C06C9C04A4B4F55DB44A0B
, sB705078CD4668BF78FEC948887DC38E7F7009BD3 : std_logic; signal s58CADDC8C7BAEBB2F1BE1E3F81F88F7A2668AC6B : std_logic := '0'; signal s7ED82462457B7203581ED9137518C167BEF13332 : std_logic_vector(1023 downto 0) := (others => '0');  signal sF3D9EE3E8A9B9537B59BF1BC9AD253A9B9B3BA6F
 : std_logic_vector(15 downto 0) := (others => '0'); signal sD002ACC5EBB2EC7EB1FC13567D61EE5BAF4CF118 : std_logic_vector( 9 downto 0) := (others => '0'); signal s2F3E7D44955F57475B683D067234C302BA0AD368 : std_logic_vector(15 downto 0) := (others => '0'); 
signal s3094B769D050989FA6EAD7EBC720891B215FA368 : std_logic_vector( 9 downto 0) := (others => '0'); signal s851F6427F4B10553861E8D231E289C621601C2B3 : std_logic_vector(15 downto 0) := (others => '0'); begin version_o <= "10" & s731A256AA7EC109FE962BF102445534C5772925D
 & s7EC4167F3F7F1E99D074313BF18FF4BA05E7ED10 & s5907A17D8E29C7EB61D4F347241BFE4DAC407AEA;  sB3DEBC4A1333AD928E577F918D84173520930691 : process(clk_i) begin if rising_edge(clk_i) then  s39BBA73E802D1EC6F9481E64A0C553405F91F14A(1) <= i_serial_clk; for s22E10B4A27DF5837B1EF92698C744643B209134E
 in 1 to s39BBA73E802D1EC6F9481E64A0C553405F91F14A'LENGTH-1 loop s39BBA73E802D1EC6F9481E64A0C553405F91F14A(s22E10B4A27DF5837B1EF92698C744643B209134E+1) <= s39BBA73E802D1EC6F9481E64A0C553405F91F14A(s22E10B4A27DF5837B1EF92698C744643B209134E); end loop; end 
if; end process sB3DEBC4A1333AD928E577F918D84173520930691;  s1BACD241F56E4F52722832FA830845B2068BC767 <= not s39BBA73E802D1EC6F9481E64A0C553405F91F14A(3) and s39BBA73E802D1EC6F9481E64A0C553405F91F14A(2); s03C86E6A8EC0C1604AE1C69CEB6A81B140CF163E <= s39BBA73E802D1EC6F9481E64A0C553405F91F14A
(3) and not s39BBA73E802D1EC6F9481E64A0C553405F91F14A(2);  sC205E4933A5E47EF50DA2E1B76E65C772A99BD19 : process(clk_i) begin if rising_edge(clk_i) then  sDD66F717A56E6D482292350AFE88447E9E2FB37F(1) <= i_serial; for s22E10B4A27DF5837B1EF92698C744643B209134E
 in 1 to sDD66F717A56E6D482292350AFE88447E9E2FB37F'LENGTH-1 loop sDD66F717A56E6D482292350AFE88447E9E2FB37F(s22E10B4A27DF5837B1EF92698C744643B209134E+1) <= sDD66F717A56E6D482292350AFE88447E9E2FB37F(s22E10B4A27DF5837B1EF92698C744643B209134E); end loop;  if 
s1BACD241F56E4F52722832FA830845B2068BC767 = '1' then s5C9DDF5B777BD5A3F655299884019D187CEB0736 <= sDD66F717A56E6D482292350AFE88447E9E2FB37F(2); end if; end if; end process sC205E4933A5E47EF50DA2E1B76E65C772A99BD19;  s5195EFEEEF3FA327D997E7C77C21627F37E4F83C
 <= sDD66F717A56E6D482292350AFE88447E9E2FB37F(2) and not s5C9DDF5B777BD5A3F655299884019D187CEB0736 and s1BACD241F56E4F52722832FA830845B2068BC767;    s20295094C230D54A994AE88B87B9386DA31BB10B : process(clk_i) begin if rising_edge(clk_i) then if reset_i='1' 
then s7437C738E80B44EBF7CA42B918E6968B6656249F <= s4EEF46B8032D06418C2A950FC6E48D5A56D77264; else s7437C738E80B44EBF7CA42B918E6968B6656249F <= s5FDA25AB9BF862813FA68F7621B5928C66206883; end if; end if; end process s20295094C230D54A994AE88B87B9386DA31BB10B
;  sE176EF29DBBED9187A59C427BC4A15DE8B881084 : process(s7437C738E80B44EBF7CA42B918E6968B6656249F, s03C86E6A8EC0C1604AE1C69CEB6A81B140CF163E, s1BACD241F56E4F52722832FA830845B2068BC767, s5195EFEEEF3FA327D997E7C77C21627F37E4F83C, s3E66115776824191EC46FFEDCE8964F683B11326
, sAABA4D54E9D1D3E0E35625A7E9DAF3FECB7C633F, s440318DC9344B28FB76FFB67D03C27AF3B02548D, sBCFB815ECFC1ADE1DD3A8C00366D0325652CDF68, tm_i, tR_i) begin  s5FDA25AB9BF862813FA68F7621B5928C66206883 <= s7437C738E80B44EBF7CA42B918E6968B6656249F;  case s7437C738E80B44EBF7CA42B918E6968B6656249F
 is  when s4EEF46B8032D06418C2A950FC6E48D5A56D77264 => if s03C86E6A8EC0C1604AE1C69CEB6A81B140CF163E = '1' then s5FDA25AB9BF862813FA68F7621B5928C66206883 <= sBB12D33790A5D3018B4D986F4ADB83977C5D8601; end if;  when sBB12D33790A5D3018B4D986F4ADB83977C5D8601 =>
 if s3E66115776824191EC46FFEDCE8964F683B11326 >= sC74718EA1B32E1BE7F9362F1CB8194555A8B7321 then s5FDA25AB9BF862813FA68F7621B5928C66206883 <= s39392447A31070974A90414173657878F7BACB37; end if;  when s39392447A31070974A90414173657878F7BACB37 => if s3E66115776824191EC46FFEDCE8964F683B11326
 >= sC1671CA18999DFAA45150AF19CC9FCDC05B45FC2 then  if s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = sB64238E7DDBD6F205572B1E9360AE1265D8B4AEA or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s577F58458D046FA77A685C62ED8B8FEF8CDC09C9 or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E
 = s552E31DD6EF995EED1A8B6C12E49DC2C0A51F02F or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = sFD1F530F2A18F9FF75CACE3E3D4051529EEF6982 or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s4BAA4FCE531A4298A40EF2ED066D556B6C1ECA42 or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E
 = sC8DFB6E167EC00F6006ED436F19C33DEA279EBB8 then s5FDA25AB9BF862813FA68F7621B5928C66206883 <= s80DC381C4925691B4334DD614AE199EF1D448C52;  else s5FDA25AB9BF862813FA68F7621B5928C66206883 <= sED64C84C9A97C77A28959EB3D8FD87CFD05499E0; end if; end if;  when s80DC381C4925691B4334DD614AE199EF1D448C52
 => if s3E66115776824191EC46FFEDCE8964F683B11326 >= s73B96A69A181F16E9161FFCBBB71691BE5986214 then s5FDA25AB9BF862813FA68F7621B5928C66206883 <= s67E7CF8001D8C888E6037A63B2A88D9E50C20BF3; end if;  when s67E7CF8001D8C888E6037A63B2A88D9E50C20BF3 => if s3E66115776824191EC46FFEDCE8964F683B11326
 >= s0C8BF396CD56CBB5C916487998FFF3E0646F0DA8 then s5FDA25AB9BF862813FA68F7621B5928C66206883 <= sED64C84C9A97C77A28959EB3D8FD87CFD05499E0; end if;  when sED64C84C9A97C77A28959EB3D8FD87CFD05499E0 => if s3E66115776824191EC46FFEDCE8964F683B11326 >= sAC85A76D3768A4693698919CFE1AC38E3EC7E60B
 then s5FDA25AB9BF862813FA68F7621B5928C66206883 <= sC8D8E0168DF0925533D8199135EDFCE49E855CE9; end if;  when sC8D8E0168DF0925533D8199135EDFCE49E855CE9 => if s440318DC9344B28FB76FFB67D03C27AF3B02548D = '1' then s5FDA25AB9BF862813FA68F7621B5928C66206883 <= s58B24B948EA83C487DAFFEC05D93C39626E147FF
; end if;  when s58B24B948EA83C487DAFFEC05D93C39626E147FF => if s3E66115776824191EC46FFEDCE8964F683B11326 >= sAABA4D54E9D1D3E0E35625A7E9DAF3FECB7C633F then  if s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s6DF2D092E032E7162C3A0DCC2D5A97E7D64555CC or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E
 = s7C44A19C549366606448A233C29ACDE5E6A81157 or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s57B57A47070F7BCB8EEBBEEA644F26DD6561AA10 or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s1BBF2B23FDB75A9E9E9C8410C6BD529018F0523E or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E
 = sEF8743F14736EEC37C81CB3F1D2B016A785A0472 or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s467E7002675271D0D9C72D30C95CAD20E650A403 then if sF74B9451531F47DEF952886360EE46EDA03FABA6 /= s83F243E9AEA0950EEEE87EEFF9FF2B8AA0412294 then s5FDA25AB9BF862813FA68F7621B5928C66206883
 <= s9361618BB4D0D11E48353A207CDF79F17E90ECC6;  elsif s10C1DD445A18FDB20BE62ADD7A9A8635E879AD33 /= s57E60BF34E25CCC564142C57DBFF63876615DB5E then s5FDA25AB9BF862813FA68F7621B5928C66206883 <= sC9891EDB20266FE6D4FB2432877D93C6F27E651B;  elsif s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E
 = s6DF2D092E032E7162C3A0DCC2D5A97E7D64555CC then s5FDA25AB9BF862813FA68F7621B5928C66206883 <= s88BB3E464A5433B5E70C481850CFB4250671F723;  else s5FDA25AB9BF862813FA68F7621B5928C66206883 <= sD1A28D5936291214869D8F06C0ADAF373A1B02C6;  end if;  else s5FDA25AB9BF862813FA68F7621B5928C66206883
 <= s88BB3E464A5433B5E70C481850CFB4250671F723;  end if; end if;  when s9361618BB4D0D11E48353A207CDF79F17E90ECC6 => if s3E66115776824191EC46FFEDCE8964F683B11326 >= sE417F33BECFBA77833DA36525F430E5AEB7C96D5 then if s10C1DD445A18FDB20BE62ADD7A9A8635E879AD33 /= 
s57E60BF34E25CCC564142C57DBFF63876615DB5E then s5FDA25AB9BF862813FA68F7621B5928C66206883 <= sC9891EDB20266FE6D4FB2432877D93C6F27E651B;  elsif s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s6DF2D092E032E7162C3A0DCC2D5A97E7D64555CC then s5FDA25AB9BF862813FA68F7621B5928C66206883
 <= s88BB3E464A5433B5E70C481850CFB4250671F723;  else s5FDA25AB9BF862813FA68F7621B5928C66206883 <= sD1A28D5936291214869D8F06C0ADAF373A1B02C6;  end if; end if;  when sC9891EDB20266FE6D4FB2432877D93C6F27E651B => if s3E66115776824191EC46FFEDCE8964F683B11326 >= 
sE417F33BECFBA77833DA36525F430E5AEB7C96D5 then if s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s6DF2D092E032E7162C3A0DCC2D5A97E7D64555CC then s5FDA25AB9BF862813FA68F7621B5928C66206883 <= s88BB3E464A5433B5E70C481850CFB4250671F723;  else s5FDA25AB9BF862813FA68F7621B5928C66206883
 <= sD1A28D5936291214869D8F06C0ADAF373A1B02C6;  end if; end if;  when sD1A28D5936291214869D8F06C0ADAF373A1B02C6 => if s3E66115776824191EC46FFEDCE8964F683B11326 >= sAC85A76D3768A4693698919CFE1AC38E3EC7E60B then s5FDA25AB9BF862813FA68F7621B5928C66206883 <= 
s1375AEE1631E1F16F7F548230C9A174D991B8343; end if;  when s1375AEE1631E1F16F7F548230C9A174D991B8343 => if s5195EFEEEF3FA327D997E7C77C21627F37E4F83C = '1' then s5FDA25AB9BF862813FA68F7621B5928C66206883 <= s51B97BD443CF4AC466F639B508697B38106C2BA3; end if;  
when s51B97BD443CF4AC466F639B508697B38106C2BA3 => if s3E66115776824191EC46FFEDCE8964F683B11326 >= s73B96A69A181F16E9161FFCBBB71691BE5986214 then s5FDA25AB9BF862813FA68F7621B5928C66206883 <= s46DB2160F9823D6161D8CD94822C414FA337C670; end if;  when s46DB2160F9823D6161D8CD94822C414FA337C670
 => if s3E66115776824191EC46FFEDCE8964F683B11326 >= s0C8BF396CD56CBB5C916487998FFF3E0646F0DA8 then s5FDA25AB9BF862813FA68F7621B5928C66206883 <= sE39C1BB78C737B4D4A9AEC7FAE586981C1DD6B52; end if;  when sE39C1BB78C737B4D4A9AEC7FAE586981C1DD6B52 => if s3E66115776824191EC46FFEDCE8964F683B11326
 >= sAC85A76D3768A4693698919CFE1AC38E3EC7E60B then s5FDA25AB9BF862813FA68F7621B5928C66206883 <= s13CF374CF3BFFB5D28DC3FA96C2EDB6E5F3847E9; end if;  when s88BB3E464A5433B5E70C481850CFB4250671F723 => if s1BACD241F56E4F52722832FA830845B2068BC767 = '1' then s5FDA25AB9BF862813FA68F7621B5928C66206883
 <= s13CF374CF3BFFB5D28DC3FA96C2EDB6E5F3847E9; end if;  when s13CF374CF3BFFB5D28DC3FA96C2EDB6E5F3847E9 => if sBCFB815ECFC1ADE1DD3A8C00366D0325652CDF68 >= unsigned(tm_i) then s5FDA25AB9BF862813FA68F7621B5928C66206883 <= sB75F5ECEEDFEADF68941469BEA18B3230DC55E12
; end if;  if s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s1E05517C0679F267FA88812F99D44A02FF4ED0F5 then if s1BACD241F56E4F52722832FA830845B2068BC767 = '1' then s5FDA25AB9BF862813FA68F7621B5928C66206883 <= sC8D8E0168DF0925533D8199135EDFCE49E855CE9; end if
; end if;  when sB75F5ECEEDFEADF68941469BEA18B3230DC55E12 => if sBCFB815ECFC1ADE1DD3A8C00366D0325652CDF68 >= unsigned(tR_i) then s5FDA25AB9BF862813FA68F7621B5928C66206883 <= s4EEF46B8032D06418C2A950FC6E48D5A56D77264; end if; when others => s5FDA25AB9BF862813FA68F7621B5928C66206883
 <= s4EEF46B8032D06418C2A950FC6E48D5A56D77264; end case;  if sBCFB815ECFC1ADE1DD3A8C00366D0325652CDF68 >= s768F8BF346D525F17E3ACF7560EB0D135C6F4041 then s5FDA25AB9BF862813FA68F7621B5928C66206883 <= s4EEF46B8032D06418C2A950FC6E48D5A56D77264; end if; end process
 sE176EF29DBBED9187A59C427BC4A15DE8B881084;   sB91AFC40BC30F66F8C035D36F1449EC546A40CF9 : process(clk_i) begin if rising_edge(clk_i) then if s1BACD241F56E4F52722832FA830845B2068BC767 = '1' then  if s7437C738E80B44EBF7CA42B918E6968B6656249F = s39392447A31070974A90414173657878F7BACB37
 then s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E <= s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E(s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E'HIGH-1 downto 0) & sDD66F717A56E6D482292350AFE88447E9E2FB37F(2); end if;   if s7437C738E80B44EBF7CA42B918E6968B6656249F = 
s80DC381C4925691B4334DD614AE199EF1D448C52 or s7437C738E80B44EBF7CA42B918E6968B6656249F = s51B97BD443CF4AC466F639B508697B38106C2BA3 then sD379CAE4835BBA8234DDEC3E02227FC8A456159E <= sD379CAE4835BBA8234DDEC3E02227FC8A456159E(sD379CAE4835BBA8234DDEC3E02227FC8A456159E
'HIGH-1 downto 0) & sDD66F717A56E6D482292350AFE88447E9E2FB37F(2); end if;   if s7437C738E80B44EBF7CA42B918E6968B6656249F = s67E7CF8001D8C888E6037A63B2A88D9E50C20BF3 or s7437C738E80B44EBF7CA42B918E6968B6656249F = s46DB2160F9823D6161D8CD94822C414FA337C670 then
 sCDC84BF1C2EA12755C5188D514BC2D52B0FD0981 <= sCDC84BF1C2EA12755C5188D514BC2D52B0FD0981(sCDC84BF1C2EA12755C5188D514BC2D52B0FD0981'HIGH-1 downto 0) & sDD66F717A56E6D482292350AFE88447E9E2FB37F(2); end if; end if; end if; end process sB91AFC40BC30F66F8C035D36F1449EC546A40CF9
;   s6B0540852F85AEF1567805B6B5FBA3EB514B1FDA : process(clk_i) begin if rising_edge(clk_i) then  if s7437C738E80B44EBF7CA42B918E6968B6656249F = sED64C84C9A97C77A28959EB3D8FD87CFD05499E0 and s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = sB64238E7DDBD6F205572B1E9360AE1265D8B4AEA
 then if sD379CAE4835BBA8234DDEC3E02227FC8A456159E(7) = '1' then s74479D486ED1C3DA5D4D8F982E552DE6F4019633 <= sD379CAE4835BBA8234DDEC3E02227FC8A456159E; end if; end if;  if s7437C738E80B44EBF7CA42B918E6968B6656249F = s46DB2160F9823D6161D8CD94822C414FA337C670
 and s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s7C44A19C549366606448A233C29ACDE5E6A81157 then if sD379CAE4835BBA8234DDEC3E02227FC8A456159E(7) = '1' then  s74479D486ED1C3DA5D4D8F982E552DE6F4019633 <= sD379CAE4835BBA8234DDEC3E02227FC8A456159E; s49778255829DFE971575864AE71D03CF1A0C4867
 <= sCDC84BF1C2EA12755C5188D514BC2D52B0FD0981(7 downto 0); else  if sD379CAE4835BBA8234DDEC3E02227FC8A456159E(7 downto 4) = X"4" then s10C1DD445A18FDB20BE62ADD7A9A8635E879AD33 <= sD379CAE4835BBA8234DDEC3E02227FC8A456159E; elsif sD379CAE4835BBA8234DDEC3E02227FC8A456159E
(7 downto 4) = X"5" then sF74B9451531F47DEF952886360EE46EDA03FABA6 <= sD379CAE4835BBA8234DDEC3E02227FC8A456159E; end if; end if; end if; end if; end process s6B0540852F85AEF1567805B6B5FBA3EB514B1FDA;    sFF8FC730077EC55526DE85F408923A3080B52842 : process(
clk_i) begin if rising_edge(clk_i) then if reset_i='1' then s1E02444D182262D00D4A327664194E0E7C9BCD58 <= s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C; else s1E02444D182262D00D4A327664194E0E7C9BCD58 <= s61E8DE0133C8A0EA7C46D3E5F1005799218FEF8B; end if; end if
; end process sFF8FC730077EC55526DE85F408923A3080B52842;  sDEE32D457486E9BDB246C33FFA400B49A7163158 : process(s1E02444D182262D00D4A327664194E0E7C9BCD58, s7437C738E80B44EBF7CA42B918E6968B6656249F, s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E, sFF8DA13899BDB1FC1B166E7DBE024EA19D9D8E78
, sFD38B58449B1F8FD27CEFABE026072920D7C6664) begin  s61E8DE0133C8A0EA7C46D3E5F1005799218FEF8B <= s1E02444D182262D00D4A327664194E0E7C9BCD58; s440318DC9344B28FB76FFB67D03C27AF3B02548D <= '0'; sF4A7A88B0CE794196EC3287991182494C4CF68BB <= '0'; case s1E02444D182262D00D4A327664194E0E7C9BCD58
 is  when s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C => if s7437C738E80B44EBF7CA42B918E6968B6656249F = sBB12D33790A5D3018B4D986F4ADB83977C5D8601 then  s61E8DE0133C8A0EA7C46D3E5F1005799218FEF8B <= s89180489BEBF665610DC5098AB8F99C0BBF612FE; end if; if s7437C738E80B44EBF7CA42B918E6968B6656249F
 = sC8D8E0168DF0925533D8199135EDFCE49E855CE9 then  sF4A7A88B0CE794196EC3287991182494C4CF68BB <= '1'; s61E8DE0133C8A0EA7C46D3E5F1005799218FEF8B <= sB72BA5545AAD812117645A3F42558C3927D9E971; end if;   when s89180489BEBF665610DC5098AB8F99C0BBF612FE => if s7437C738E80B44EBF7CA42B918E6968B6656249F
 = sED64C84C9A97C77A28959EB3D8FD87CFD05499E0 then  if s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = sB64238E7DDBD6F205572B1E9360AE1265D8B4AEA or  s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s4BAA4FCE531A4298A40EF2ED066D556B6C1ECA42 then  sF4A7A88B0CE794196EC3287991182494C4CF68BB
 <= '1';  s61E8DE0133C8A0EA7C46D3E5F1005799218FEF8B <= sF0D99209603F6F7473DE58A048ABB74800BF9B6E; else s61E8DE0133C8A0EA7C46D3E5F1005799218FEF8B <= sE73FCB3053E16A73428686A101357781139D2C9D;  end if; end if;  when sF0D99209603F6F7473DE58A048ABB74800BF9B6E
 => if sFF8DA13899BDB1FC1B166E7DBE024EA19D9D8E78 >= s7F754F692527BC0267C69BBEFF22B0EB623D725D then s61E8DE0133C8A0EA7C46D3E5F1005799218FEF8B <= s0FC3DA9494BAFC3ED1F299DDF23029966E219F55; end if;  when sB72BA5545AAD812117645A3F42558C3927D9E971 => if sFF8DA13899BDB1FC1B166E7DBE024EA19D9D8E78
 >= s180C3B3A658D0B94ADDD3EBA8B3FD02288454264 then s61E8DE0133C8A0EA7C46D3E5F1005799218FEF8B <= s0FC3DA9494BAFC3ED1F299DDF23029966E219F55; end if;  when sE73FCB3053E16A73428686A101357781139D2C9D => if sFD38B58449B1F8FD27CEFABE026072920D7C6664 >= s8A2992E6D362DBB70C96CD6B71F48399524E30D2
 then s61E8DE0133C8A0EA7C46D3E5F1005799218FEF8B <= s0FC3DA9494BAFC3ED1F299DDF23029966E219F55; end if;  when s0FC3DA9494BAFC3ED1F299DDF23029966E219F55 => s440318DC9344B28FB76FFB67D03C27AF3B02548D <= '1'; if s7437C738E80B44EBF7CA42B918E6968B6656249F = s58B24B948EA83C487DAFFEC05D93C39626E147FF
 then s61E8DE0133C8A0EA7C46D3E5F1005799218FEF8B <= s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C; end if; when others => s61E8DE0133C8A0EA7C46D3E5F1005799218FEF8B <= s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C; end case; end process sDEE32D457486E9BDB246C33FFA400B49A7163158
;   sFD179360A8EF07805D297F2F18EDD591576A6974 : process(clk_i) begin if rising_edge(clk_i) then   if to_integer(signed(sFF8DA13899BDB1FC1B166E7DBE024EA19D9D8E78)) /= -1 then if s1BACD241F56E4F52722832FA830845B2068BC767 = '1' then sFF8DA13899BDB1FC1B166E7DBE024EA19D9D8E78
 <= sFF8DA13899BDB1FC1B166E7DBE024EA19D9D8E78 + 1; end if; end if;  if sF4A7A88B0CE794196EC3287991182494C4CF68BB = '1' then sFF8DA13899BDB1FC1B166E7DBE024EA19D9D8E78 <= (others => '0'); end if;   if to_integer(signed(sFD38B58449B1F8FD27CEFABE026072920D7C6664
)) /= -1 then sFD38B58449B1F8FD27CEFABE026072920D7C6664 <= sFD38B58449B1F8FD27CEFABE026072920D7C6664 + 1; end if;  if s7437C738E80B44EBF7CA42B918E6968B6656249F /= sBB12D33790A5D3018B4D986F4ADB83977C5D8601 and s5FDA25AB9BF862813FA68F7621B5928C66206883 = sBB12D33790A5D3018B4D986F4ADB83977C5D8601
 then sFD38B58449B1F8FD27CEFABE026072920D7C6664 <= (others => '0'); end if;   if s7437C738E80B44EBF7CA42B918E6968B6656249F = sED64C84C9A97C77A28959EB3D8FD87CFD05499E0 then s8A2992E6D362DBB70C96CD6B71F48399524E30D2 <= unsigned(tcal_i(21 downto 0));  if s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E
 = s552E31DD6EF995EED1A8B6C12E49DC2C0A51F02F or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s577F58458D046FA77A685C62ED8B8FEF8CDC09C9 or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = sC8DFB6E167EC00F6006ED436F19C33DEA279EBB8 then  s8A2992E6D362DBB70C96CD6B71F48399524E30D2
 <= sB6C4B6996BE4000D3F7E6A44BB9ED1B6A592CAF0; end if; if s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = sFD1F530F2A18F9FF75CACE3E3D4051529EEF6982 then  s8A2992E6D362DBB70C96CD6B71F48399524E30D2 <= sD0F92C1D45611463356A15CFF87B99280A8A24F1; end if; end if;  
 if to_integer(signed(s3E66115776824191EC46FFEDCE8964F683B11326)) /= -1 then if s1BACD241F56E4F52722832FA830845B2068BC767 = '1' then s3E66115776824191EC46FFEDCE8964F683B11326 <= s3E66115776824191EC46FFEDCE8964F683B11326 + 1; end if; end if;  if s7437C738E80B44EBF7CA42B918E6968B6656249F
 /= s5FDA25AB9BF862813FA68F7621B5928C66206883 then s3E66115776824191EC46FFEDCE8964F683B11326 <= (others => '0'); end if;   if to_integer(signed(sBCFB815ECFC1ADE1DD3A8C00366D0325652CDF68)) /= -1 then sBCFB815ECFC1ADE1DD3A8C00366D0325652CDF68 <= sBCFB815ECFC1ADE1DD3A8C00366D0325652CDF68
 + 1; end if;  if s7437C738E80B44EBF7CA42B918E6968B6656249F /= s5FDA25AB9BF862813FA68F7621B5928C66206883 or s7437C738E80B44EBF7CA42B918E6968B6656249F = s4EEF46B8032D06418C2A950FC6E48D5A56D77264 then sBCFB815ECFC1ADE1DD3A8C00366D0325652CDF68 <= (others => '0');
 end if;  if s7437C738E80B44EBF7CA42B918E6968B6656249F /= s4EEF46B8032D06418C2A950FC6E48D5A56D77264 and s5FDA25AB9BF862813FA68F7621B5928C66206883 = s4EEF46B8032D06418C2A950FC6E48D5A56D77264 then s34682EDE73B453730FDDB73AE693BF6858792888 <= s34682EDE73B453730FDDB73AE693BF6858792888
 + 1; end if; end if; end process sFD179360A8EF07805D297F2F18EDD591576A6974;    s0399AD38FFE6E9911310CCF2C7975E26207D5D3D <= to_integer(unsigned(numPulPosVal_i));    sAABA4D54E9D1D3E0E35625A7E9DAF3FECB7C633F <= to_unsigned(30, 6) when s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E
 = sB64238E7DDBD6F205572B1E9360AE1265D8B4AEA or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s552E31DD6EF995EED1A8B6C12E49DC2C0A51F02F or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s577F58458D046FA77A685C62ED8B8FEF8CDC09C9 or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E
 = sFD1F530F2A18F9FF75CACE3E3D4051529EEF6982 or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s4BAA4FCE531A4298A40EF2ED066D556B6C1ECA42 or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = sC8DFB6E167EC00F6006ED436F19C33DEA279EBB8 else  to_unsigned(2 + s0399AD38FFE6E9911310CCF2C7975E26207D5D3D
 + 5, 6) when s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s1E05517C0679F267FA88812F99D44A02FF4ED0F5 else  to_unsigned(3 + s0399AD38FFE6E9911310CCF2C7975E26207D5D3D + 5, 6) when s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s6DF2D092E032E7162C3A0DCC2D5A97E7D64555CC
 or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s7C44A19C549366606448A233C29ACDE5E6A81157 or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s57B57A47070F7BCB8EEBBEEA644F26DD6561AA10 or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s1BBF2B23FDB75A9E9E9C8410C6BD529018F0523E
 or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = sEF8743F14736EEC37C81CB3F1D2B016A785A0472 or s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E = s467E7002675271D0D9C72D30C95CAD20E650A403 else  to_unsigned(1 + 40 + 5, 6) when s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E
 = s1E05517C0679F267FA88812F99D44A02FF4ED0F5 else  (others => '0');  sD2575E546E2EC143C5C4DD4FCD988505DC92A552 <= dataRx_MSB_i(15 downto 0) & dataRx_LSB_i(31 downto 0); sCFD226CC0ECDD9D07EE7E693ABB8A3A3B1E2CF73(47 downto 16) <= (others => '0') when dataMode_i
(0) = '1' else sD2575E546E2EC143C5C4DD4FCD988505DC92A552(47 downto 16); sCFD226CC0ECDD9D07EE7E693ABB8A3A3B1E2CF73(15 downto 0) <= std_logic_vector(s34682EDE73B453730FDDB73AE693BF6858792888) when dataMode_i(0) = '1' else sD2575E546E2EC143C5C4DD4FCD988505DC92A552
(15 downto 0);  s06D292C2A3FDB9DCE32D576C2C85F8ED0E615CE9: for s5C5D67AB466573ED99CC2706B41FF2D01C569AAD in sCFD226CC0ECDD9D07EE7E693ABB8A3A3B1E2CF73'range generate sEE8C5684D6E32E443D201C83D1FDFBBBAC150FAD(sEE8C5684D6E32E443D201C83D1FDFBBBAC150FAD'HIGH - 
s5C5D67AB466573ED99CC2706B41FF2D01C569AAD) <= sCFD226CC0ECDD9D07EE7E693ABB8A3A3B1E2CF73(s5C5D67AB466573ED99CC2706B41FF2D01C569AAD); end generate;  sC4B6EA407C3AA8DD2E6A18E7F77C14FACC951414 <= dataMode_i(2); s06E676C0BDF7C68FD7495790A14A2FEBA13D3DB6 <= dataMode_i
(3); warning <= dataMode_i(4); s76804DD01BB29A387010BCE68256FDB2A4020735 <= '1'; sCB42C2FDABBD75F13A77BB4E139059E0A23744FD <= '0';  sD98C8E6D4E6D4476AF57C3F9E1684609B34E6FB7 : process(s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E, sD379CAE4835BBA8234DDEC3E02227FC8A456159E
, sC4B6EA407C3AA8DD2E6A18E7F77C14FACC951414, s06E676C0BDF7C68FD7495790A14A2FEBA13D3DB6, sEE8C5684D6E32E443D201C83D1FDFBBBAC150FAD, s0399AD38FFE6E9911310CCF2C7975E26207D5D3D, sF3D9EE3E8A9B9537B59BF1BC9AD253A9B9B3BA6F, sCDC84BF1C2EA12755C5188D514BC2D52B0FD0981
) begin  sBB999F79F35F7555095A7373986DE0689DE5FC46 <= (others => '0'); sBB999F79F35F7555095A7373986DE0689DE5FC46(50) <= sED14BC4B3908B6DB77B3D546FFC4257CF3675A4F; case s7285EAB431F245D6C89C51D95316E4DE4AEDFC3E is  when s1E05517C0679F267FA88812F99D44A02FF4ED0F5
 => sBB999F79F35F7555095A7373986DE0689DE5FC46(49) <= sC4B6EA407C3AA8DD2E6A18E7F77C14FACC951414; sBB999F79F35F7555095A7373986DE0689DE5FC46(48 downto 1) <= sEE8C5684D6E32E443D201C83D1FDFBBBAC150FAD;  when s6DF2D092E032E7162C3A0DCC2D5A97E7D64555CC | s7C44A19C549366606448A233C29ACDE5E6A81157
 | s57B57A47070F7BCB8EEBBEEA644F26DD6561AA10 | s1BBF2B23FDB75A9E9E9C8410C6BD529018F0523E | sEF8743F14736EEC37C81CB3F1D2B016A785A0472 | s467E7002675271D0D9C72D30C95CAD20E650A403 => sBB999F79F35F7555095A7373986DE0689DE5FC46(49) <= sC4B6EA407C3AA8DD2E6A18E7F77C14FACC951414
; sBB999F79F35F7555095A7373986DE0689DE5FC46(48) <= not s06E676C0BDF7C68FD7495790A14A2FEBA13D3DB6; sBB999F79F35F7555095A7373986DE0689DE5FC46(47 downto 0) <= sEE8C5684D6E32E443D201C83D1FDFBBBAC150FAD;  when sB64238E7DDBD6F205572B1E9360AE1265D8B4AEA | s577F58458D046FA77A685C62ED8B8FEF8CDC09C9
 | sFD1F530F2A18F9FF75CACE3E3D4051529EEF6982 | s4BAA4FCE531A4298A40EF2ED066D556B6C1ECA42 | sC8DFB6E167EC00F6006ED436F19C33DEA279EBB8 => sBB999F79F35F7555095A7373986DE0689DE5FC46(49 downto 26) <= sD379CAE4835BBA8234DDEC3E02227FC8A456159E & sCDC84BF1C2EA12755C5188D514BC2D52B0FD0981
;  when s552E31DD6EF995EED1A8B6C12E49DC2C0A51F02F => sBB999F79F35F7555095A7373986DE0689DE5FC46(49 downto 26) <= sD379CAE4835BBA8234DDEC3E02227FC8A456159E & sF3D9EE3E8A9B9537B59BF1BC9AD253A9B9B3BA6F;  when s3CE74FA91201742DE9903A95D23643FE5849757A => sBB999F79F35F7555095A7373986DE0689DE5FC46
(49 downto 9) <= sC4B6EA407C3AA8DD2E6A18E7F77C14FACC951414 & X"123456789A";  when others => sBB999F79F35F7555095A7373986DE0689DE5FC46(50 downto 0) <= (others => '0'); end case; end process sD98C8E6D4E6D4476AF57C3F9E1684609B34E6FB7;  sDEBE07749EE39C0C6AE751A310A9B1432D4FAB77
 : process(s10C1DD445A18FDB20BE62ADD7A9A8635E879AD33, sD379CAE4835BBA8234DDEC3E02227FC8A456159E, warning, s76804DD01BB29A387010BCE68256FDB2A4020735, sCB42C2FDABBD75F13A77BB4E139059E0A23744FD, sF3D9EE3E8A9B9537B59BF1BC9AD253A9B9B3BA6F, s74479D486ED1C3DA5D4D8F982E552DE6F4019633
) begin  sEF80C7392E78A56484621A1127C5B6AB5F281091 <= (others => '0'); sEF80C7392E78A56484621A1127C5B6AB5F281091(24) <= not sED14BC4B3908B6DB77B3D546FFC4257CF3675A4F; sEF80C7392E78A56484621A1127C5B6AB5F281091(23) <= warning; sEF80C7392E78A56484621A1127C5B6AB5F281091
(22) <= s76804DD01BB29A387010BCE68256FDB2A4020735; sEF80C7392E78A56484621A1127C5B6AB5F281091(21) <= sCB42C2FDABBD75F13A77BB4E139059E0A23744FD; sEF80C7392E78A56484621A1127C5B6AB5F281091(20 downto 16) <= s10C1DD445A18FDB20BE62ADD7A9A8635E879AD33(4 downto 0);
 case s10C1DD445A18FDB20BE62ADD7A9A8635E879AD33 is when sC467071B4163DF3B730A3D8FDBA24B62A24337A7 => sEF80C7392E78A56484621A1127C5B6AB5F281091(15 downto 0) <= X"0000"; when s497A41403D0E1204014E9B612AD737C8D35B3826 => sEF80C7392E78A56484621A1127C5B6AB5F281091
(15 downto 0) <= X"0000"; when sFA0C0FC5DB4F0920FD931E78C8F3FFB13715D3FD => sEF80C7392E78A56484621A1127C5B6AB5F281091(15 downto 0) <= X"0011"; when s0E620B5ED6FCC4C01B20B593ADCB3709FA0BE26E => sEF80C7392E78A56484621A1127C5B6AB5F281091(15 downto 0) <= X"0110";
 when s5AE40AED79A09E5B98B32D981F056406C9D6D977 => sEF80C7392E78A56484621A1127C5B6AB5F281091(15 downto 0) <= X"1100"; when sF76D4DB16EF1ADE5770C213F52561503D34DEF48 => sEF80C7392E78A56484621A1127C5B6AB5F281091(15 downto 0) <= sD379CAE4835BBA8234DDEC3E02227FC8A456159E
 & sF3D9EE3E8A9B9537B59BF1BC9AD253A9B9B3BA6F(7 downto 0); when sFE54C7D0CC6A2E8CFA4216501DCE1D8F436FEDC6 => sEF80C7392E78A56484621A1127C5B6AB5F281091(15 downto 0) <= sD379CAE4835BBA8234DDEC3E02227FC8A456159E & sF3D9EE3E8A9B9537B59BF1BC9AD253A9B9B3BA6F(15 
downto 8); when s7840E41D30357FC6180671D694922360D68CC896 => sEF80C7392E78A56484621A1127C5B6AB5F281091(15 downto 0) <= sD379CAE4835BBA8234DDEC3E02227FC8A456159E & s74479D486ED1C3DA5D4D8F982E552DE6F4019633; when sB8FBD8D6BBEDF46E31A0507EABC8F686CFB5CFA0 => 
sEF80C7392E78A56484621A1127C5B6AB5F281091(15 downto 0) <= sD379CAE4835BBA8234DDEC3E02227FC8A456159E & X"FE"; when s41500258240C5111284D79C684750BDFCF9BB4C9 => sEF80C7392E78A56484621A1127C5B6AB5F281091(15 downto 0) <= X"0022"; when s726B1776BF9E9357377F4BD979D5C542A12D7ECE
 => sEF80C7392E78A56484621A1127C5B6AB5F281091(15 downto 0) <= X"0220"; when s83ADFBE2A97ACC106909DAC843AFC39378B31F29 => sEF80C7392E78A56484621A1127C5B6AB5F281091(15 downto 0) <= X"2200"; when sCF680DC8F214E3DEE1C42E950A30559BBAC4F3EB => sEF80C7392E78A56484621A1127C5B6AB5F281091
(15 downto 0) <= temperature_i(15 downto 0); when s030F867793634A136982960F35AEAEFADF3FF2E0 => sEF80C7392E78A56484621A1127C5B6AB5F281091(15 downto 0) <= temperature_i(15 downto 0); when sDB159321904E6E9F130985F9B9AA585A8C6A0047 => sEF80C7392E78A56484621A1127C5B6AB5F281091
(15 downto 0) <= X"AD5E"; when s57E60BF34E25CCC564142C57DBFF63876615DB5E => sEF80C7392E78A56484621A1127C5B6AB5F281091(15 downto 0) <= X"EE33"; when others => sEF80C7392E78A56484621A1127C5B6AB5F281091(15 downto 0) <= (others => '0'); end case; end process 
sDEBE07749EE39C0C6AE751A310A9B1432D4FAB77;  s3F3D358D7C358CDDAD537D0CCCB2CA2150153B9A : process(sF74B9451531F47DEF952886360EE46EDA03FABA6, warning, s76804DD01BB29A387010BCE68256FDB2A4020735, sCB42C2FDABBD75F13A77BB4E139059E0A23744FD) begin  sDDFA38A34F7901FE6E261DE887A8F537753CF545
 <= (others => '0'); sDDFA38A34F7901FE6E261DE887A8F537753CF545(24) <= not sED14BC4B3908B6DB77B3D546FFC4257CF3675A4F; sDDFA38A34F7901FE6E261DE887A8F537753CF545(23) <= warning; sDDFA38A34F7901FE6E261DE887A8F537753CF545(22) <= s76804DD01BB29A387010BCE68256FDB2A4020735
; sDDFA38A34F7901FE6E261DE887A8F537753CF545(21) <= sCB42C2FDABBD75F13A77BB4E139059E0A23744FD; sDDFA38A34F7901FE6E261DE887A8F537753CF545(20 downto 16) <= sF74B9451531F47DEF952886360EE46EDA03FABA6(4 downto 0); case sF74B9451531F47DEF952886360EE46EDA03FABA6 
is when s190163C428AF25FC3187CA8FA8195F66129DEE18 => sDDFA38A34F7901FE6E261DE887A8F537753CF545(15 downto 0) <= X"0000"; when sD753454CEAEA82A91076ECB6EF4A5F2112BC34A0 => sDDFA38A34F7901FE6E261DE887A8F537753CF545(15 downto 0) <= commutation_i(7 downto 0) & x"00";
 when sF99D1A97BFDA9B5076280F23CECAAF884FCBA996 => sDDFA38A34F7901FE6E261DE887A8F537753CF545(15 downto 0) <= X"0011"; when s51302044F211B9E83B0E4160532E89D41D26179F => sDDFA38A34F7901FE6E261DE887A8F537753CF545(15 downto 0) <= commutation_i(7 downto 0) & x"11";
 when sA0E09E1DFA0715EA5072265E84B3B90BDEF4A330 => sDDFA38A34F7901FE6E261DE887A8F537753CF545(15 downto 0) <= X"C000"; when s98D7FC4F26467AB3B384D5297B7DAA0066EAB130 => sDDFA38A34F7901FE6E261DE887A8F537753CF545(15 downto 0) <= X"C011"; when s57A7C76B0F0C0E6103B6BDE4922267DFC1C6CAC8
 => sDDFA38A34F7901FE6E261DE887A8F537753CF545(15 downto 0) <= X"0022"; when sFAEE7C7664BC579F00801F34E53AA70BD65A7874 => sDDFA38A34F7901FE6E261DE887A8F537753CF545(15 downto 0) <= X"0220"; when s1E153525FB86CE60222E8A7CBAA485AF861B1D74 => sDDFA38A34F7901FE6E261DE887A8F537753CF545
(15 downto 0) <= X"2200"; when s27FC1A1F329912801D6E9215F3007A63A8623499 => sDDFA38A34F7901FE6E261DE887A8F537753CF545(15 downto 0) <= X"0000"; when sE312DD9AD97739BDE32B25BD07E6F495A41E9C6F => sDDFA38A34F7901FE6E261DE887A8F537753CF545(15 downto 0) <= X"AFFE";
 when s97161BEE2D29B3E48064B3B437D9507452C8BE43 => sDDFA38A34F7901FE6E261DE887A8F537753CF545(15 downto 0) <= X"B00B"; when s83F243E9AEA0950EEEE87EEFF9FF2B8AA0412294 => sDDFA38A34F7901FE6E261DE887A8F537753CF545(15 downto 0) <= X"C0DE"; when others => sDDFA38A34F7901FE6E261DE887A8F537753CF545
(15 downto 0) <= (others => '0'); end case; end process s3F3D358D7C358CDDAD537D0CCCB2CA2150153B9A;  sB705078CD4668BF78FEC948887DC38E7F7009BD3 <= ((s63B7F7C57F075889730F3ADD94597ABD229977FB(4) and sD3C21919EB55E97996C06C9C04A4B4F55DB44A0B) xor sAE11F5A23788CBD8FAF306A52CAC70458125557A
(50)) when s7437C738E80B44EBF7CA42B918E6968B6656249F = s58B24B948EA83C487DAFFEC05D93C39626E147FF else ((s63B7F7C57F075889730F3ADD94597ABD229977FB(4) and sD3C21919EB55E97996C06C9C04A4B4F55DB44A0B) xor sCFF2D518C744D824B9DE2B4D9AFBF5F4725457B2(24)) when s7437C738E80B44EBF7CA42B918E6968B6656249F
 = sC9891EDB20266FE6D4FB2432877D93C6F27E651B else ((s63B7F7C57F075889730F3ADD94597ABD229977FB(4) and sD3C21919EB55E97996C06C9C04A4B4F55DB44A0B) xor sB355DE414F49CCFFF6381B960907D94AA7FBF024(24)) when s7437C738E80B44EBF7CA42B918E6968B6656249F = s9361618BB4D0D11E48353A207CDF79F17E90ECC6
 else '0'; sD3C21919EB55E97996C06C9C04A4B4F55DB44A0B <= '1';   sD1A14F957B86B32C91CEFE47296C70BA09C866F7 : process(clk_i) begin if rising_edge(clk_i) then  if s7437C738E80B44EBF7CA42B918E6968B6656249F = sC8D8E0168DF0925533D8199135EDFCE49E855CE9 then sAE11F5A23788CBD8FAF306A52CAC70458125557A
 <= sBB999F79F35F7555095A7373986DE0689DE5FC46; sCFF2D518C744D824B9DE2B4D9AFBF5F4725457B2 <= sEF80C7392E78A56484621A1127C5B6AB5F281091; sB355DE414F49CCFFF6381B960907D94AA7FBF024 <= sDDFA38A34F7901FE6E261DE887A8F537753CF545; end if;  if s1BACD241F56E4F52722832FA830845B2068BC767
 = '1' then  if s7437C738E80B44EBF7CA42B918E6968B6656249F = s58B24B948EA83C487DAFFEC05D93C39626E147FF or s7437C738E80B44EBF7CA42B918E6968B6656249F = sC9891EDB20266FE6D4FB2432877D93C6F27E651B or s7437C738E80B44EBF7CA42B918E6968B6656249F = s9361618BB4D0D11E48353A207CDF79F17E90ECC6
 then  if (s7437C738E80B44EBF7CA42B918E6968B6656249F = s58B24B948EA83C487DAFFEC05D93C39626E147FF and (s3E66115776824191EC46FFEDCE8964F683B11326 < sAABA4D54E9D1D3E0E35625A7E9DAF3FECB7C633F-5)) or (s7437C738E80B44EBF7CA42B918E6968B6656249F /= s58B24B948EA83C487DAFFEC05D93C39626E147FF
 and (s3E66115776824191EC46FFEDCE8964F683B11326 < sE417F33BECFBA77833DA36525F430E5AEB7C96D5-5)) then  if s3E66115776824191EC46FFEDCE8964F683B11326 >= 1 then s63B7F7C57F075889730F3ADD94597ABD229977FB(4) <= s63B7F7C57F075889730F3ADD94597ABD229977FB(3); s63B7F7C57F075889730F3ADD94597ABD229977FB
(3) <= ((sB705078CD4668BF78FEC948887DC38E7F7009BD3 and sD3C21919EB55E97996C06C9C04A4B4F55DB44A0B) xor s63B7F7C57F075889730F3ADD94597ABD229977FB(2)); s63B7F7C57F075889730F3ADD94597ABD229977FB(2) <= s63B7F7C57F075889730F3ADD94597ABD229977FB(1); s63B7F7C57F075889730F3ADD94597ABD229977FB
(1) <= ((sB705078CD4668BF78FEC948887DC38E7F7009BD3 and sD3C21919EB55E97996C06C9C04A4B4F55DB44A0B) xor s63B7F7C57F075889730F3ADD94597ABD229977FB(0)); s63B7F7C57F075889730F3ADD94597ABD229977FB(0) <= sB705078CD4668BF78FEC948887DC38E7F7009BD3; end if;  if s7437C738E80B44EBF7CA42B918E6968B6656249F
 = s58B24B948EA83C487DAFFEC05D93C39626E147FF then s58CADDC8C7BAEBB2F1BE1E3F81F88F7A2668AC6B <= sAE11F5A23788CBD8FAF306A52CAC70458125557A(sAE11F5A23788CBD8FAF306A52CAC70458125557A'HIGH); sAE11F5A23788CBD8FAF306A52CAC70458125557A <= sAE11F5A23788CBD8FAF306A52CAC70458125557A
(sAE11F5A23788CBD8FAF306A52CAC70458125557A'HIGH-1 downto 0) & '0';  elsif s7437C738E80B44EBF7CA42B918E6968B6656249F = sC9891EDB20266FE6D4FB2432877D93C6F27E651B then s58CADDC8C7BAEBB2F1BE1E3F81F88F7A2668AC6B <= sCFF2D518C744D824B9DE2B4D9AFBF5F4725457B2(sCFF2D518C744D824B9DE2B4D9AFBF5F4725457B2
'HIGH); sCFF2D518C744D824B9DE2B4D9AFBF5F4725457B2 <= sCFF2D518C744D824B9DE2B4D9AFBF5F4725457B2(sCFF2D518C744D824B9DE2B4D9AFBF5F4725457B2'HIGH-1 downto 0) & '0';  else s58CADDC8C7BAEBB2F1BE1E3F81F88F7A2668AC6B <= sB355DE414F49CCFFF6381B960907D94AA7FBF024(sB355DE414F49CCFFF6381B960907D94AA7FBF024
'HIGH); sB355DE414F49CCFFF6381B960907D94AA7FBF024 <= sB355DE414F49CCFFF6381B960907D94AA7FBF024(sB355DE414F49CCFFF6381B960907D94AA7FBF024'HIGH-1 downto 0) & '0'; end if;  else s58CADDC8C7BAEBB2F1BE1E3F81F88F7A2668AC6B <= not s63B7F7C57F075889730F3ADD94597ABD229977FB
(4) xor dataMode_i(1);  s63B7F7C57F075889730F3ADD94597ABD229977FB <= s63B7F7C57F075889730F3ADD94597ABD229977FB(3 downto 0) & '1';  end if; end if;  if s7437C738E80B44EBF7CA42B918E6968B6656249F = sE39C1BB78C737B4D4A9AEC7FAE586981C1DD6B52 or s7437C738E80B44EBF7CA42B918E6968B6656249F
 = sD1A28D5936291214869D8F06C0ADAF373A1B02C6 then s58CADDC8C7BAEBB2F1BE1E3F81F88F7A2668AC6B <= '1'; end if;  if s7437C738E80B44EBF7CA42B918E6968B6656249F = s1375AEE1631E1F16F7F548230C9A174D991B8343 then s58CADDC8C7BAEBB2F1BE1E3F81F88F7A2668AC6B <= '0'; end
 if; end if;   if s7437C738E80B44EBF7CA42B918E6968B6656249F = s13CF374CF3BFFB5D28DC3FA96C2EDB6E5F3847E9 then s58CADDC8C7BAEBB2F1BE1E3F81F88F7A2668AC6B <= '1'; end if;  if s7437C738E80B44EBF7CA42B918E6968B6656249F = sB75F5ECEEDFEADF68941469BEA18B3230DC55E12
 or s7437C738E80B44EBF7CA42B918E6968B6656249F = s4EEF46B8032D06418C2A950FC6E48D5A56D77264 then s58CADDC8C7BAEBB2F1BE1E3F81F88F7A2668AC6B <= '0'; end if;    if s7437C738E80B44EBF7CA42B918E6968B6656249F = s4EEF46B8032D06418C2A950FC6E48D5A56D77264 then o_drive_en
 <= '1'; end if;  if s7437C738E80B44EBF7CA42B918E6968B6656249F=sBB12D33790A5D3018B4D986F4ADB83977C5D8601 then o_drive_en <= '0'; end if;  if s7437C738E80B44EBF7CA42B918E6968B6656249F = sED64C84C9A97C77A28959EB3D8FD87CFD05499E0 or s7437C738E80B44EBF7CA42B918E6968B6656249F
 = sE39C1BB78C737B4D4A9AEC7FAE586981C1DD6B52 then if s3E66115776824191EC46FFEDCE8964F683B11326=x"00000001" then  if s03C86E6A8EC0C1604AE1C69CEB6A81B140CF163E='1' then  o_drive_en <= '1'; end if; end if; end if;  if s7437C738E80B44EBF7CA42B918E6968B6656249F
 = sD1A28D5936291214869D8F06C0ADAF373A1B02C6 then if s3E66115776824191EC46FFEDCE8964F683B11326=x"00000002" then  if s03C86E6A8EC0C1604AE1C69CEB6A81B140CF163E='1' then  o_drive_en <= '0'; end if; end if; end if; end if; end process sD1A14F957B86B32C91CEFE47296C70BA09C866F7
; s45C9B0206D487B36E381524C94D668132932FD0D: process(clk_i)  begin if rising_edge(clk_i) then  s7ED82462457B7203581ED9137518C167BEF13332 <= s7ED82462457B7203581ED9137518C167BEF13332(1022 downto 0) & s58CADDC8C7BAEBB2F1BE1E3F81F88F7A2668AC6B;   o_serial <= 
s7ED82462457B7203581ED9137518C167BEF13332(to_integer(unsigned(td_i(9 downto 0)))); end if; end process s45C9B0206D487B36E381524C94D668132932FD0D;    sF9E69889EF39BA019E2115826DF2A9EC0FCBF7CB: process(clk_i) begin if rising_edge(clk_i) then  case s74479D486ED1C3DA5D4D8F982E552DE6F4019633
 is  when X"B9" => if unsigned(sD379CAE4835BBA8234DDEC3E02227FC8A456159E) < 4 then sD002ACC5EBB2EC7EB1FC13567D61EE5BAF4CF118 <= "00000000" & sD379CAE4835BBA8234DDEC3E02227FC8A456159E(1 downto 0); end if;  when X"A1" => if unsigned(sD379CAE4835BBA8234DDEC3E02227FC8A456159E
) > 3 and unsigned(sD379CAE4835BBA8234DDEC3E02227FC8A456159E) < 16 then sD002ACC5EBB2EC7EB1FC13567D61EE5BAF4CF118 <= "000000" & sD379CAE4835BBA8234DDEC3E02227FC8A456159E(3 downto 0); end if;  when X"A3" => if unsigned(sD379CAE4835BBA8234DDEC3E02227FC8A456159E
) < 16 then sD002ACC5EBB2EC7EB1FC13567D61EE5BAF4CF118 <= "000001" & sD379CAE4835BBA8234DDEC3E02227FC8A456159E(3 downto 0); end if;  when X"A5" => if unsigned(sD379CAE4835BBA8234DDEC3E02227FC8A456159E) < 16 then sD002ACC5EBB2EC7EB1FC13567D61EE5BAF4CF118 <= "000010" & 
sD379CAE4835BBA8234DDEC3E02227FC8A456159E(3 downto 0); end if;  when X"A7" => if unsigned(sD379CAE4835BBA8234DDEC3E02227FC8A456159E) < 16 then sD002ACC5EBB2EC7EB1FC13567D61EE5BAF4CF118(5 downto 0) <= "11" & sD379CAE4835BBA8234DDEC3E02227FC8A456159E(3 downto
 0); end if;  when X"A9" => if unsigned(sD379CAE4835BBA8234DDEC3E02227FC8A456159E) > 63 then sD002ACC5EBB2EC7EB1FC13567D61EE5BAF4CF118 <= "00" & sD379CAE4835BBA8234DDEC3E02227FC8A456159E; end if;  when X"AB" => sD002ACC5EBB2EC7EB1FC13567D61EE5BAF4CF118 <= "01" & 
sD379CAE4835BBA8234DDEC3E02227FC8A456159E;  when X"AD" => sD002ACC5EBB2EC7EB1FC13567D61EE5BAF4CF118 <= "10" & sD379CAE4835BBA8234DDEC3E02227FC8A456159E;          when X"B7" => sD002ACC5EBB2EC7EB1FC13567D61EE5BAF4CF118 <= "11" & sD379CAE4835BBA8234DDEC3E02227FC8A456159E
;  when X"BD" => if unsigned(sD379CAE4835BBA8234DDEC3E02227FC8A456159E) < 63 then s3094B769D050989FA6EAD7EBC720891B215FA368 <= "00" & sD379CAE4835BBA8234DDEC3E02227FC8A456159E; end if;  when X"BB" => s3094B769D050989FA6EAD7EBC720891B215FA368 <= "01" & sD379CAE4835BBA8234DDEC3E02227FC8A456159E
;  when X"BF" => if unsigned(s49778255829DFE971575864AE71D03CF1A0C4867) < 2 then s3094B769D050989FA6EAD7EBC720891B215FA368 <= '1' & s49778255829DFE971575864AE71D03CF1A0C4867(0) & sD379CAE4835BBA8234DDEC3E02227FC8A456159E; end if; when others => NULL; end 
case s74479D486ED1C3DA5D4D8F982E552DE6F4019633;  s2F3E7D44955F57475B683D067234C302BA0AD368 <= s1CFD18110A517486D9B5DAED3C58733F8D80465E(to_integer(unsigned(sD002ACC5EBB2EC7EB1FC13567D61EE5BAF4CF118))); s851F6427F4B10553861E8D231E289C621601C2B3 <= sCD229F113F7E82913D1F47B1ED664487BEEB48A8
(to_integer(unsigned(s3094B769D050989FA6EAD7EBC720891B215FA368)));   if s74479D486ED1C3DA5D4D8F982E552DE6F4019633 = X"A1" and sD379CAE4835BBA8234DDEC3E02227FC8A456159E = X"0D" then sF3D9EE3E8A9B9537B59BF1BC9AD253A9B9B3BA6F <= '1' & numPulPosVal_i(14 downto
 0);  elsif s74479D486ED1C3DA5D4D8F982E552DE6F4019633 = X"A3" and sD379CAE4835BBA8234DDEC3E02227FC8A456159E = X"01" then sF3D9EE3E8A9B9537B59BF1BC9AD253A9B9B3BA6F <= distRev_i(15 downto 0);  elsif s74479D486ED1C3DA5D4D8F982E552DE6F4019633 = X"A7" and sD379CAE4835BBA8234DDEC3E02227FC8A456159E
 = X"0F" then sF3D9EE3E8A9B9537B59BF1BC9AD253A9B9B3BA6F <= std_logic_vector(unsigned(s2F3E7D44955F57475B683D067234C302BA0AD368) + unsigned(numPulPosVal_i(14 downto 0)) + unsigned(distRev_i(15 downto 0)));  elsif s74479D486ED1C3DA5D4D8F982E552DE6F4019633 = X"B9" 
then sF3D9EE3E8A9B9537B59BF1BC9AD253A9B9B3BA6F <= X"0000";  elsif s74479D486ED1C3DA5D4D8F982E552DE6F4019633 = X"BF" or s74479D486ED1C3DA5D4D8F982E552DE6F4019633 = X"BD" or s74479D486ED1C3DA5D4D8F982E552DE6F4019633 = X"BB" then sF3D9EE3E8A9B9537B59BF1BC9AD253A9B9B3BA6F
 <= s851F6427F4B10553861E8D231E289C621601C2B3;  else sF3D9EE3E8A9B9537B59BF1BC9AD253A9B9B3BA6F <= s2F3E7D44955F57475B683D067234C302BA0AD368; end if; end if; end process sF9E69889EF39BA019E2115826DF2A9EC0FCBF7CB; end struct; 