--*******************************************************************************************
--
--                                                          endatreduced
--                                                          ==========
-- File Name:        endatreduced.vhd
-- Project:          Endat Reduced
-- Modul Name:       ---
-- Author:           Frank Seiler/ MAZeT GmbH
--                   MAZeT GmbH
--                   Goeschwitzer Strasse 32        
--                   D-07745 Jena
--
-- Specification:    ---
--                                                             
-- Synthesis:        (Tested with Synoplfy 8.6.2) 
--                              
-- Script:           ENDAT22.prj
--                               
-- Simulation:       Cadence NCVHDL V3.41, V5.1
-- 
-- Function:         EnDat Reduced
--                                  
-- History: F.Seiler xx.12.2007 Initial Version EnDat2.1 only
--          F.Seiler xx.07.2008 AddOn EnDat2.2
--          F.Seiler 17.09.2008 some signals renamed 
--*******************************************************************************************
library ieee; use ieee.std_logic_1164.all; use ieee.std_logic_unsigned.all; USE ieee.std_logic_arith.CONV_STD_LOGIC_VECTOR; use ieee.std_logic_misc.all; use ieee.numeric_std.all; entity endatreduced is generic ( sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81 : 
integer:= 6;  s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95 : integer:= 7;  s2B661762AEA08905D55D9C993A5A3B37FF2EC6CD : integer:= 32;  sCD3268FB2E69A058B357988C1BAD31C26B18C0D3 : integer:= 56;   s4A8616F7DBB06E84D521DFE24490E8ADB037CBB1 : boolean:= false;  s745F184CD6754435326632E8F885833C3FD28CAA
 : integer:= 2);  port ( s82C78E3CD667612DE97ED7C5FA8365F21045093F : in std_logic;  sF1FC47B36F2DA843714A618883F345968A471A76 : in std_logic;   sF4DBC68D16423B9DD337E166EF77471DCEA3D993 : in std_logic;  s298D55696DC353303493AAE18ABFD0C95B97F0F7 : out std_logic
;  s858AFDE712A6913772203E81B3BDEEB1165DDD96 : out std_logic;  s1504ADD95BA0488B2CA487398BBC3A3FB56ED3A4 : out std_logic;   sAF6F101406809B45BE51F9E400AB99C6466D8AAE: in integer;  s11183BFF0C2D855AEA5F48EC192129844E5C157D: in integer;  s940FAE140F86D7AAE5446A4FA8C953A8EA6B637D
 : in integer;  sDF43AA73D6AFC95DE6173B25BC8316E2AE46E705 : in integer;  s7F693B395683971F9F003DC8983DF2304C3CE968 : in std_logic;  s90196555A8BFC1A5EE5D4925FBA2AF598F9D76F9: in std_logic_vector(1 downto 0);   sE420A02AD972A785E332BF27D04B53B8868A4F0E : in
 std_logic_vector(s2B661762AEA08905D55D9C993A5A3B37FF2EC6CD -1 downto 0);  s86F6EB29E2D65A736372F43D1F449BCF6DB2BA0A : in std_logic;  sA16C86782D377069727114AB99F123218DC1EE4E : out std_logic;  s07A72EEC7FE78460042B89F4D0DA7BE551FEC90A : out std_logic;  s28EDCB4BE5AFFD576E337FA1A3A5AAEEA7D7B33C
 : out std_logic;  s353B8D288425991916C61A5A9DFE44B11BBCF753 : out std_logic_vector(sCD3268FB2E69A058B357988C1BAD31C26B18C0D3 -1 downto 0);  s43F7D19F6FFB52EF969FC2858BC1CA57C001562A : out std_logic_vector( 4 downto 0);  sC4B6EA407C3AA8DD2E6A18E7F77C14FACC951414
 : out std_logic;  s06E676C0BDF7C68FD7495790A14A2FEBA13D3DB6 : out std_logic;  s0BFFA2AEF006C5821760F1A640F5456669E1486A : out std_logic;  s32CF03224D0C548C4F44A5420AF0E47F9CE9CB0F : out std_logic;  s601E9D380BAA3E6CC5A2AEE58C2C073DF7C885D1 : out std_logic
;  sA516DA7C751934DBE51FECC222FA4984B32B3692 : out std_logic;  s7975BCABF4261F33B14B8E6E764BC7741562D89E : out std_logic;  s7DC4BA5492A3997AE8E131EA0BD60F3CED572BBD: in std_logic;  s1B88525B5C44F4D86E63397D61F66E7B1225355E : out std_logic_vector(63 downto
 0);  s8ABB29C3748C74A80027187254C15F46F51EF2A2 : out std_logic_vector(3 downto 0);  s83F675DB784B205945DE32DEA0270B2CF41801FE : out std_logic_vector(s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95 -1 downto 0)  ); end endatreduced; Architecture s75BE5DEF24CA4A61B9676CCF1CC90EBA505DC89E
 of endatreduced is component pdm generic ( s8012194BD35F0878CACF167A77EE7A04F42ED698 : integer:= 5;  s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95 : integer:= 7;   s4A8616F7DBB06E84D521DFE24490E8ADB037CBB1 : boolean:= false;  s745F184CD6754435326632E8F885833C3FD28CAA
 : integer:= 2);  port ( s82C78E3CD667612DE97ED7C5FA8365F21045093F : in std_logic;  sF1FC47B36F2DA843714A618883F345968A471A76 : in std_logic;   sA73098C7B13AE4EE2D18DD1A3C28A605F0315F7B : in std_logic;  s90196555A8BFC1A5EE5D4925FBA2AF598F9D76F9: in std_logic_vector
(1 downto 0);  pdm : in std_logic;  sA871AC5299DD9A2B5922B93C415099F5B17A2CAA: in std_logic_vector( 3 downto 0);  s3DE9704ED5E8C46005ACD085579D848AC14D5B18 : in std_logic;  s3878B21E042F1AD8CD97DB6E7D00908A99649D03 : in std_logic;  s134B4B78A794B9AC71D2041279723343FA183008
 : in std_logic;  s264475A303AC7031FBC8591205A50743DAEAD9CA : in std_logic;  s125623D1F098599393E5DE6A762EFFC9DACED467 : out std_logic;  s3943BBC49DABABC540DBFCA8F53E255877F4D8F1 : out std_logic_vector(s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95 -1 downto 0); 
 sC95BB2A3A95288115289D986565E400E04F2B5A0 : out std_logic;  s79CBDE1F1AE76DE1CEAD5B67EFDA2C6953987F5C: out std_logic; sEA5E54196582D991021F5AB19DAC58C70947FB22: out std_logic_vector(s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95 -1 downto 0); s1B88525B5C44F4D86E63397D61F66E7B1225355E
 : out std_logic_vector(63 downto 0);   s11183BFF0C2D855AEA5F48EC192129844E5C157D: in integer;  s940FAE140F86D7AAE5446A4FA8C953A8EA6B637D : in integer  ); end component; signal sA871AC5299DD9A2B5922B93C415099F5B17A2CAA: std_logic_vector( 3 downto 0); signal
 s0C95BB05F974B637452566ABF145558806623663, s90FD026CDBD878ABC461660ADF31E80BA177A2AA, s6A18EECF6FABFF8383A93194D7C565C57343844A: std_logic; signal s67A0998548ED967361FBF09931BE2B937104D248, s49807CD868D22833D34695DE61B3DA5F68DD41DC: std_logic; signal sCBF7A0249B3E467C859DC6110B4A5C709856666B
, sA8F3D27EFD5141F07A5CE1B87DA29A4ABD9AF24E, s69B82088412476FAF1B1D1362493AAF169716766: std_logic; signal sDE7CDC6FDA2463F07579EEEE09153F29DF743435, s776F81CD2516996DEA92F16B486A7FED89C09EB8, sA03ED9A8ADD1D6369CFFD09A3B204681F4FD4323: std_logic; signal s92A8540F7FAAFAFEC21E720F4DA706442BB74A1F
,s1D698942AE29B843C12FC388FE7AE002990CA8DC,s7B2460199CAF56FF7F3235463ED56BE379DEF304: std_logic; signal s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9: std_logic_vector(sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81 -1 downto 0); signal sDE3723024059B3D9CCBE053F62FD7805FEF750D5
: std_logic_vector(s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95 -1 downto 0); signal s3DE9704ED5E8C46005ACD085579D848AC14D5B18, s8DB4E21FE7FB3394A51B5A83BE1F618408AEC221: std_logic; signal sC5B8A229B10A712ADBC43679D961A8B4B2922490 : std_logic; signal s69C5A9568767AD2BF8234062710212C330AC69A1
 : std_logic; signal s3878B21E042F1AD8CD97DB6E7D00908A99649D03: std_logic; signal s73124B1BDDFA8E0A4B7A0970B215A0C89FD997AA: std_logic; signal s8949CFA6A16FC99FBD129BE88F26A12A41A2ACE1: std_logic; signal sD24BF1A9310E03CA3B5DBECC807B894C04E87F42: std_logic
; signal s5995FA7F6E2087033AB6935283687FAE3F27CA76: std_logic; signal sCBB4558CFEFE324102C5417B1E5A0CBDB858B168, sCAF301BC43AEA5B1C0FCEBF9360CAC2EDDDEF3D5: std_logic_vector(sCD3268FB2E69A058B357988C1BAD31C26B18C0D3 downto 0); signal s06C5EFDBF86E27179DFD37C48A46E20937862C9D
: std_logic_vector(sCD3268FB2E69A058B357988C1BAD31C26B18C0D3 +1 downto 0); signal s1792FD2BB24BFB0793974D92FA74B345EB0CCAF3 : std_logic; signal s064596695B62E7458EDC8A508E0EE076015E8499, s2324B84C04CC4C838C23EB219AAB9CF288E9F546: std_logic; signal s01BC98CC8DA65101EC29BFBE486670F7247144FB
 : std_logic; signal sBC134FF3B7F8A030502858E6E7D1EF2141E3647D: std_logic; signal sFCFAEC304D530FD8874F63BC093FFA6D2F2C9E57: std_logic_vector(s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95 -1 downto 0); signal s566CCC14B9C50B000C4DB011CD7D548338128B26: std_logic_vector
(s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95 -1 downto 0); signal sE9B685CB6A496C918D983B7EC72C8D3D8EC3123B : std_logic; signal s264475A303AC7031FBC8591205A50743DAEAD9CA: std_logic_vector(3 downto 0); signal s48925532037BE5F8C053A6D5DB7767BB7A703DCF: std_logic
; signal s46B3B4D75B1901ADCD5C39F1B58D398BB213B6BF: std_logic; signal s134B4B78A794B9AC71D2041279723343FA183008: std_logic; signal s035B34BD1D4E71D6E05E7E0C12748A22F2AB0BAF: std_logic; signal s7A68704BA3FEDFAA8EBAC048D2067E5B0158325F: std_logic_vector(sCD3268FB2E69A058B357988C1BAD31C26B18C0D3
 -1 downto 0); signal s0572647003D0AE885FEB3E9760C0F5C78BA6B52A: integer; signal sB2FF42C79B0D014AFEDA0B7415287448CC5F1553: integer; signal s1FAAEBEE7B845D3CBACD553CA078AD4D43E0ADFA, sC1AA6E43EDA79EA468391A422C8C0A84CAFE4DD9: std_logic; signal s4045C346006E7236123346044B3C0BBE00D1391F
: std_logic; signal s27D6EF4CA3309F1B892E6207A8D14DCC6F949466: std_logic; signal s63DCD945122E83C803DEB91867786995FFCFE62A: std_logic; signal s78D1CF9FDB871B9B4256DCE09B67D406079A5FB8: std_logic; signal s9606968BB22D6E6CABE7FC03219FFECDA4CB919D, s228AB3A49C983930DA44D78299DB703391BE79F3
: std_logic_vector( 4 downto 0); signal s74009442A8C13802B71EA10AB67B2A147A944F36: std_logic_vector( 4 downto 0); signal s3C3AD1732E30E3202F031BD11ADED227CB12BDB6: std_logic_vector( 4 downto 0);  signal sD3C21919EB55E97996C06C9C04A4B4F55DB44A0B, s8507177FCFDBD094828F65353CFC1170B6FEA614
: std_logic; signal s3751FAFD204DD6237D01F1ABA4489435D55D9525: std_logic; signal sC280108DF6F82A156D03BC60D309452D917A55B9: std_logic_vector(s745F184CD6754435326632E8F885833C3FD28CAA -1 downto 0); signal sAEF369739F02576F7BA2574212961A3126F4E307, s54A764BE0E3DFF5AFCCB0617D1E670FDF5B430FC
: std_logic; signal s6A5FE1CD0E944495E6BF7242D05EAEACFBA89ACF, s125623D1F098599393E5DE6A762EFFC9DACED467: std_logic; signal sBE3694D6DE3020DED7EF579482C5628CB0A7D85D, s9279E19351BBF8CD9801F2005A998BF5C72988B9 : std_logic; signal sAA4741C86EC7F1A9388F089FDAFF07D1332CA196
: std_logic; signal sE734111027AE4A3C909A98A63E7589D18CBEA161: std_logic_vector(s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95 -1 downto 0); signal s01AF22A3811BAB6264C575A96A22B593A64576AE, s425754F7414052216602B6E7EA8CE966DBE28995: std_logic; signal s3943BBC49DABABC540DBFCA8F53E255877F4D8F1
: std_logic_vector(s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95 -1 downto 0); signal sC95BB2A3A95288115289D986565E400E04F2B5A0 : std_logic;  signal s013E9FFBF04A31B71784E98EAB7A683996BA039E : std_logic_vector(sCD3268FB2E69A058B357988C1BAD31C26B18C0D3 -1 downto
 0); signal s03384791D53DA7C796CA8B60E2BF84B83EF294E1, s34D0BA0417C5C46CBC3249708B1E4BB573BE4F13 : std_logic; signal s3FE6E74D86F2DF0268B67C717D22E60D521CE7E5, s3B95BCD02DFA6D86D669FA75993367A9B3D3207A : std_logic; signal sD02015CB26E1B7025DF2F7880CFEB9376D504E69
, s855750D5D93589BB5ABD95DCDECD97BED3D7389E : std_logic; signal sEA8188CAD31707F17B299650F81C67D601FE09D7 : std_logic_vector(5 downto 0); signal sA73098C7B13AE4EE2D18DD1A3C28A605F0315F7B : std_logic; begin s7A68704BA3FEDFAA8EBAC048D2067E5B0158325F <= CONV_STD_LOGIC_VECTOR
(0, sCD3268FB2E69A058B357988C1BAD31C26B18C0D3); s6A5FE1CD0E944495E6BF7242D05EAEACFBA89ACF <= s7F693B395683971F9F003DC8983DF2304C3CE968;  process(s82C78E3CD667612DE97ED7C5FA8365F21045093F) begin if rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then
 if sF1FC47B36F2DA843714A618883F345968A471A76 = '0' then s5995FA7F6E2087033AB6935283687FAE3F27CA76 <= '0'; else case sA871AC5299DD9A2B5922B93C415099F5B17A2CAA is when "0000" => if s86F6EB29E2D65A736372F43D1F449BCF6DB2BA0A = '1' then s5995FA7F6E2087033AB6935283687FAE3F27CA76
 <= '1'; end if; when "1111" => s5995FA7F6E2087033AB6935283687FAE3F27CA76 <= '0'; when others => s5995FA7F6E2087033AB6935283687FAE3F27CA76 <= s5995FA7F6E2087033AB6935283687FAE3F27CA76; end case; end if; end if; end process;  process(s82C78E3CD667612DE97ED7C5FA8365F21045093F
) begin if rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then if sF1FC47B36F2DA843714A618883F345968A471A76 = '0' then sA871AC5299DD9A2B5922B93C415099F5B17A2CAA <= "0000"; s49807CD868D22833D34695DE61B3DA5F68DD41DC <= '0'; s69B82088412476FAF1B1D1362493AAF169716766
 <= '0'; sA03ED9A8ADD1D6369CFFD09A3B204681F4FD4323 <= '0'; s7B2460199CAF56FF7F3235463ED56BE379DEF304 <= '0'; sA8F3D27EFD5141F07A5CE1B87DA29A4ABD9AF24E <= '0'; s776F81CD2516996DEA92F16B486A7FED89C09EB8 <= '0'; s1D698942AE29B843C12FC388FE7AE002990CA8DC <= '0'; else s49807CD868D22833D34695DE61B3DA5F68DD41DC <= s67A0998548ED967361FBF09931BE2B937104D248; s69B82088412476FAF1B1D1362493AAF169716766 <= sA8F3D27EFD5141F07A5CE1B87DA29A4ABD9AF24E; sA03ED9A8ADD1D6369CFFD09A3B204681F4FD4323 <= s776F81CD2516996DEA92F16B486A7FED89C09EB8
; s7B2460199CAF56FF7F3235463ED56BE379DEF304 <= s1D698942AE29B843C12FC388FE7AE002990CA8DC; sA8F3D27EFD5141F07A5CE1B87DA29A4ABD9AF24E <= sCBF7A0249B3E467C859DC6110B4A5C709856666B; s776F81CD2516996DEA92F16B486A7FED89C09EB8 <= sDE7CDC6FDA2463F07579EEEE09153F29DF743435
; s1D698942AE29B843C12FC388FE7AE002990CA8DC <= s92A8540F7FAAFAFEC21E720F4DA706442BB74A1F; case sA871AC5299DD9A2B5922B93C415099F5B17A2CAA is when "0000" =>  if s8DB4E21FE7FB3394A51B5A83BE1F618408AEC221 = '1' and s5995FA7F6E2087033AB6935283687FAE3F27CA76 = '1' 
then sA871AC5299DD9A2B5922B93C415099F5B17A2CAA <= "0001"; end if; when "0001" =>  if s3878B21E042F1AD8CD97DB6E7D00908A99649D03 = '0' then if sC5B8A229B10A712ADBC43679D961A8B4B2922490 = '1' then if s8DB4E21FE7FB3394A51B5A83BE1F618408AEC221 = '1' then sA871AC5299DD9A2B5922B93C415099F5B17A2CAA
 <= "0010"; end if; end if; end if; when "0010" | "0100" | "1010" | "1011" | "1101" | "1110" =>  if s3878B21E042F1AD8CD97DB6E7D00908A99649D03 = '0' then if sC5B8A229B10A712ADBC43679D961A8B4B2922490 = '1' then if s8DB4E21FE7FB3394A51B5A83BE1F618408AEC221 = '1' 
then sA871AC5299DD9A2B5922B93C415099F5B17A2CAA <= sA871AC5299DD9A2B5922B93C415099F5B17A2CAA + '1'; end if; end if; end if; when "0011" =>  if s3878B21E042F1AD8CD97DB6E7D00908A99649D03 = '1' then if sC5B8A229B10A712ADBC43679D961A8B4B2922490 = '1' then if s8DB4E21FE7FB3394A51B5A83BE1F618408AEC221
 = '1' then sA871AC5299DD9A2B5922B93C415099F5B17A2CAA <= sA871AC5299DD9A2B5922B93C415099F5B17A2CAA + '1'; end if; end if; end if; when "0101" =>  if s125623D1F098599393E5DE6A762EFFC9DACED467 = '0' or s6A5FE1CD0E944495E6BF7242D05EAEACFBA89ACF = '0' then if
 s3878B21E042F1AD8CD97DB6E7D00908A99649D03 = '0' then if sC5B8A229B10A712ADBC43679D961A8B4B2922490 = '1' then if s8DB4E21FE7FB3394A51B5A83BE1F618408AEC221 = '1' then if s90196555A8BFC1A5EE5D4925FBA2AF598F9D76F9 /= "00" then sA871AC5299DD9A2B5922B93C415099F5B17A2CAA
 <= "1000"; else if sA73098C7B13AE4EE2D18DD1A3C28A605F0315F7B = '0' then sA871AC5299DD9A2B5922B93C415099F5B17A2CAA <= "1111";  else sA871AC5299DD9A2B5922B93C415099F5B17A2CAA <= "1010";  end if; end if; end if; end if; end if; end if; if s125623D1F098599393E5DE6A762EFFC9DACED467
 = '1' and s6A5FE1CD0E944495E6BF7242D05EAEACFBA89ACF ='1' then if sAA4741C86EC7F1A9388F089FDAFF07D1332CA196 = '1' then  if sC5B8A229B10A712ADBC43679D961A8B4B2922490 = '1' then if s425754F7414052216602B6E7EA8CE966DBE28995 = '1' then  if s90196555A8BFC1A5EE5D4925FBA2AF598F9D76F9
 /= "00" then sA871AC5299DD9A2B5922B93C415099F5B17A2CAA <= "1000"; else if sA73098C7B13AE4EE2D18DD1A3C28A605F0315F7B = '0' then sA871AC5299DD9A2B5922B93C415099F5B17A2CAA <= "1111";  else sA871AC5299DD9A2B5922B93C415099F5B17A2CAA <= "1010";  end if; end if
; end if; end if; end if; end if; when "1000" =>  if s3878B21E042F1AD8CD97DB6E7D00908A99649D03 = '0' then if sC5B8A229B10A712ADBC43679D961A8B4B2922490 = '1' then if s8DB4E21FE7FB3394A51B5A83BE1F618408AEC221 = '1' then if s90196555A8BFC1A5EE5D4925FBA2AF598F9D76F9
 = "10" then sA871AC5299DD9A2B5922B93C415099F5B17A2CAA <= "1001"; else if sA73098C7B13AE4EE2D18DD1A3C28A605F0315F7B = '0' then sA871AC5299DD9A2B5922B93C415099F5B17A2CAA <= "1111";  else sA871AC5299DD9A2B5922B93C415099F5B17A2CAA <= "1010";  end if; end if; end if; end if; end if; when "1001" =>  if s3878B21E042F1AD8CD97DB6E7D00908A99649D03 = '0' then if sC5B8A229B10A712ADBC43679D961A8B4B2922490 = '1' then if s8DB4E21FE7FB3394A51B5A83BE1F618408AEC221 = '1' then if sA73098C7B13AE4EE2D18DD1A3C28A605F0315F7B = '0' 
then sA871AC5299DD9A2B5922B93C415099F5B17A2CAA <= "1111";  else sA871AC5299DD9A2B5922B93C415099F5B17A2CAA <= "1010";  end if; end if; end if; end if; when "1100" =>  if s3878B21E042F1AD8CD97DB6E7D00908A99649D03 = '0' then if sC5B8A229B10A712ADBC43679D961A8B4B2922490
 = '1' then if s8DB4E21FE7FB3394A51B5A83BE1F618408AEC221 = '1' then sA871AC5299DD9A2B5922B93C415099F5B17A2CAA <= "1101"; end if; end if; end if; when others => sA871AC5299DD9A2B5922B93C415099F5B17A2CAA <= "0000"; end case; end if; end if; end process; s0C95BB05F974B637452566ABF145558806623663
 <= '1' when sA871AC5299DD9A2B5922B93C415099F5B17A2CAA = "0001" else '0'; s67A0998548ED967361FBF09931BE2B937104D248 <= '1' when sA871AC5299DD9A2B5922B93C415099F5B17A2CAA = "0101" else '0'; sCBF7A0249B3E467C859DC6110B4A5C709856666B <= '1' when sA871AC5299DD9A2B5922B93C415099F5B17A2CAA
 = "1000" else '0'; sDE7CDC6FDA2463F07579EEEE09153F29DF743435 <= '1' when sA871AC5299DD9A2B5922B93C415099F5B17A2CAA = "1001" else '0'; s6A18EECF6FABFF8383A93194D7C565C57343844A <= '1' when sA871AC5299DD9A2B5922B93C415099F5B17A2CAA = "1100" else '0'; s92A8540F7FAAFAFEC21E720F4DA706442BB74A1F
 <= '1' when sA871AC5299DD9A2B5922B93C415099F5B17A2CAA = "1010" else '0'; s90FD026CDBD878ABC461660ADF31E80BA177A2AA <= '1' when sA871AC5299DD9A2B5922B93C415099F5B17A2CAA = "1011" else '0';   process(s82C78E3CD667612DE97ED7C5FA8365F21045093F) begin if rising_edge
(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then if sF1FC47B36F2DA843714A618883F345968A471A76 = '0' then s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 <= (others=>'0'); sD24BF1A9310E03CA3B5DBECC807B894C04E87F42 <= '0'; else if s5995FA7F6E2087033AB6935283687FAE3F27CA76
 = '1' then if s3878B21E042F1AD8CD97DB6E7D00908A99649D03 = '0' then if s3DE9704ED5E8C46005ACD085579D848AC14D5B18 = '1' then case sA871AC5299DD9A2B5922B93C415099F5B17A2CAA is when "0000" => s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 <= CONV_STD_LOGIC_VECTOR
(sAF6F101406809B45BE51F9E400AB99C6466D8AAE,sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81);  sD24BF1A9310E03CA3B5DBECC807B894C04E87F42 <= '0';  when "0001" =>  if s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 = CONV_STD_LOGIC_VECTOR(0, sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81
) then s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 <= CONV_STD_LOGIC_VECTOR(sAF6F101406809B45BE51F9E400AB99C6466D8AAE,sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81);  sD24BF1A9310E03CA3B5DBECC807B894C04E87F42 <= '1'; else s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9
 <= s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 - '1'; end if; when "0010" => sD24BF1A9310E03CA3B5DBECC807B894C04E87F42 <= '0';  when "0101" =>  if s125623D1F098599393E5DE6A762EFFC9DACED467 = '0' or s6A5FE1CD0E944495E6BF7242D05EAEACFBA89ACF = '0' then if s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9
 = CONV_STD_LOGIC_VECTOR(0, sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81) then s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 <= CONV_STD_LOGIC_VECTOR(s11183BFF0C2D855AEA5F48EC192129844E5C157D,sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81);  elsif s134B4B78A794B9AC71D2041279723343FA183008
 = '1' or s48925532037BE5F8C053A6D5DB7767BB7A703DCF = '1' then s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 <= s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 - '1'; end if; end if;  when "1000" | "1001" =>  if s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 = CONV_STD_LOGIC_VECTOR
( 0, sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81) then s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 <= CONV_STD_LOGIC_VECTOR(29, sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81);  elsif s134B4B78A794B9AC71D2041279723343FA183008 = '1' or s48925532037BE5F8C053A6D5DB7767BB7A703DCF
 = '1' then s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 <= s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 - '1'; end if;  when "1100" =>  if s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 = CONV_STD_LOGIC_VECTOR(0, sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81) then s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9
 <= CONV_STD_LOGIC_VECTOR(27,sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81);  sD24BF1A9310E03CA3B5DBECC807B894C04E87F42 <= '1'; else s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 <= s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 - '1'; sD24BF1A9310E03CA3B5DBECC807B894C04E87F42
 <= '1'; end if; when "1110" => sD24BF1A9310E03CA3B5DBECC807B894C04E87F42 <= '0';  when others => s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 <= CONV_STD_LOGIC_VECTOR(0,sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81);  end case; end if; end if; if s125623D1F098599393E5DE6A762EFFC9DACED467
 = '1' and s6A5FE1CD0E944495E6BF7242D05EAEACFBA89ACF ='1' then if sA871AC5299DD9A2B5922B93C415099F5B17A2CAA = "0101" then if sAA4741C86EC7F1A9388F089FDAFF07D1332CA196 = '1' then if s01AF22A3811BAB6264C575A96A22B593A64576AE = '1' then  if s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9
 = CONV_STD_LOGIC_VECTOR(0, sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81) then s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 <= CONV_STD_LOGIC_VECTOR(s11183BFF0C2D855AEA5F48EC192129844E5C157D,sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81);  elsif s134B4B78A794B9AC71D2041279723343FA183008
 = '1' or s48925532037BE5F8C053A6D5DB7767BB7A703DCF = '1' then s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 <= s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 - '1'; end if; end if; end if; end if; end if; end if; end if; end if; end process; sC5B8A229B10A712ADBC43679D961A8B4B2922490
 <= '1' when s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 = CONV_STD_LOGIC_VECTOR (0, sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81) else '0';   process(s82C78E3CD667612DE97ED7C5FA8365F21045093F) begin if rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then
 if sF1FC47B36F2DA843714A618883F345968A471A76 = '0' then sDE3723024059B3D9CCBE053F62FD7805FEF750D5 <= (others=>'0'); else if s1FAAEBEE7B845D3CBACD553CA078AD4D43E0ADFA = '1' and s92A8540F7FAAFAFEC21E720F4DA706442BB74A1F = '0' then sDE3723024059B3D9CCBE053F62FD7805FEF750D5
 <= (others=>'0'); elsif s86F6EB29E2D65A736372F43D1F449BCF6DB2BA0A = '1' or s5995FA7F6E2087033AB6935283687FAE3F27CA76 = '0' then  sDE3723024059B3D9CCBE053F62FD7805FEF750D5 <= CONV_STD_LOGIC_VECTOR(s0572647003D0AE885FEB3E9760C0F5C78BA6B52A, s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95
);  elsif s86F6EB29E2D65A736372F43D1F449BCF6DB2BA0A = '1' or s5995FA7F6E2087033AB6935283687FAE3F27CA76 = '1' then if sDE3723024059B3D9CCBE053F62FD7805FEF750D5 = CONV_STD_LOGIC_VECTOR(0, s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95) then sDE3723024059B3D9CCBE053F62FD7805FEF750D5
 <= CONV_STD_LOGIC_VECTOR(s0572647003D0AE885FEB3E9760C0F5C78BA6B52A, s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95);  else sDE3723024059B3D9CCBE053F62FD7805FEF750D5 <= sDE3723024059B3D9CCBE053F62FD7805FEF750D5 - '1'; end if; end if; end if; end if; end process
; sB2FF42C79B0D014AFEDA0B7415287448CC5F1553 <= sDF43AA73D6AFC95DE6173B25BC8316E2AE46E705 when s125623D1F098599393E5DE6A762EFFC9DACED467 = '0' else to_integer(unsigned(s3943BBC49DABABC540DBFCA8F53E255877F4D8F1)); s0572647003D0AE885FEB3E9760C0F5C78BA6B52A <= 
sB2FF42C79B0D014AFEDA0B7415287448CC5F1553 when sA871AC5299DD9A2B5922B93C415099F5B17A2CAA = "0000" else  sB2FF42C79B0D014AFEDA0B7415287448CC5F1553 when sA871AC5299DD9A2B5922B93C415099F5B17A2CAA = "0100" else  s940FAE140F86D7AAE5446A4FA8C953A8EA6B637D - 1; 
 s3DE9704ED5E8C46005ACD085579D848AC14D5B18 <= '1' when sDE3723024059B3D9CCBE053F62FD7805FEF750D5 = CONV_STD_LOGIC_VECTOR (0, s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95) else '0'; s8DB4E21FE7FB3394A51B5A83BE1F618408AEC221 <= '1' when sDE3723024059B3D9CCBE053F62FD7805FEF750D5
 = CONV_STD_LOGIC_VECTOR (1, s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95) else '0';  s01AF22A3811BAB6264C575A96A22B593A64576AE <= '1' when sE734111027AE4A3C909A98A63E7589D18CBEA161 = CONV_STD_LOGIC_VECTOR (0, s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95) else '0'; 
s425754F7414052216602B6E7EA8CE966DBE28995 <= '1' when sE734111027AE4A3C909A98A63E7589D18CBEA161 = CONV_STD_LOGIC_VECTOR (1, s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95) else '0';   process(s82C78E3CD667612DE97ED7C5FA8365F21045093F) begin if rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F
) then if sF1FC47B36F2DA843714A618883F345968A471A76 = '0' then s3878B21E042F1AD8CD97DB6E7D00908A99649D03 <= '1'; s73124B1BDDFA8E0A4B7A0970B215A0C89FD997AA <= '1'; else case sA871AC5299DD9A2B5922B93C415099F5B17A2CAA is when "0000" => if s86F6EB29E2D65A736372F43D1F449BCF6DB2BA0A
 = '1' then s3878B21E042F1AD8CD97DB6E7D00908A99649D03 <= '0'; s73124B1BDDFA8E0A4B7A0970B215A0C89FD997AA <= '0'; end if; when others => if s5995FA7F6E2087033AB6935283687FAE3F27CA76 = '1' then if s3DE9704ED5E8C46005ACD085579D848AC14D5B18 = '1' then s3878B21E042F1AD8CD97DB6E7D00908A99649D03
 <= not s3878B21E042F1AD8CD97DB6E7D00908A99649D03; end if; if s3DE9704ED5E8C46005ACD085579D848AC14D5B18 = '1' and sC95BB2A3A95288115289D986565E400E04F2B5A0 = '0' then s73124B1BDDFA8E0A4B7A0970B215A0C89FD997AA <= not s73124B1BDDFA8E0A4B7A0970B215A0C89FD997AA
; end if; end if; end case; end if; end if; end process;   s925915C161CC45CDD933AFAC5B654D2AD743161B: for s020F5125771EEEB6F963720A8BB968FCA977AA41 in sCBB4558CFEFE324102C5417B1E5A0CBDB858B168'range generate s29849470D152FDE2CAF8EEAB3FF07395D472D891: process
(s11183BFF0C2D855AEA5F48EC192129844E5C157D, sCBB4558CFEFE324102C5417B1E5A0CBDB858B168, sF4DBC68D16423B9DD337E166EF77471DCEA3D993) begin if s020F5125771EEEB6F963720A8BB968FCA977AA41 < (s11183BFF0C2D855AEA5F48EC192129844E5C157D) then sCAF301BC43AEA5B1C0FCEBF9360CAC2EDDDEF3D5
(s020F5125771EEEB6F963720A8BB968FCA977AA41) <= sCBB4558CFEFE324102C5417B1E5A0CBDB858B168(s020F5125771EEEB6F963720A8BB968FCA977AA41); elsif s020F5125771EEEB6F963720A8BB968FCA977AA41 = (s11183BFF0C2D855AEA5F48EC192129844E5C157D) then sCAF301BC43AEA5B1C0FCEBF9360CAC2EDDDEF3D5
(s020F5125771EEEB6F963720A8BB968FCA977AA41) <= sF4DBC68D16423B9DD337E166EF77471DCEA3D993; else sCAF301BC43AEA5B1C0FCEBF9360CAC2EDDDEF3D5(s020F5125771EEEB6F963720A8BB968FCA977AA41) <= '0'; end if; end process s29849470D152FDE2CAF8EEAB3FF07395D472D891; end 
generate;  process(s82C78E3CD667612DE97ED7C5FA8365F21045093F) begin if rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then if sF1FC47B36F2DA843714A618883F345968A471A76 = '0' then sCBB4558CFEFE324102C5417B1E5A0CBDB858B168 <= (others=>'0'); s01BC98CC8DA65101EC29BFBE486670F7247144FB
 <= '0'; s3C3AD1732E30E3202F031BD11ADED227CB12BDB6 <= (others=>'0') ; else s01BC98CC8DA65101EC29BFBE486670F7247144FB <= s064596695B62E7458EDC8A508E0EE076015E8499; if s5995FA7F6E2087033AB6935283687FAE3F27CA76 = '0' and s86F6EB29E2D65A736372F43D1F449BCF6DB2BA0A
 = '1' then sCBB4558CFEFE324102C5417B1E5A0CBDB858B168 <= '0' & sE420A02AD972A785E332BF27D04B53B8868A4F0E(s2B661762AEA08905D55D9C993A5A3B37FF2EC6CD -1 downto 0) & s7A68704BA3FEDFAA8EBAC048D2067E5B0158325F(sCD3268FB2E69A058B357988C1BAD31C26B18C0D3 - s2B661762AEA08905D55D9C993A5A3B37FF2EC6CD
 -1 downto 0);  end if; if s90FD026CDBD878ABC461660ADF31E80BA177A2AA = '1' then sCBB4558CFEFE324102C5417B1E5A0CBDB858B168 <= '0' & sE420A02AD972A785E332BF27D04B53B8868A4F0E(s2B661762AEA08905D55D9C993A5A3B37FF2EC6CD -1 downto 0) & s7A68704BA3FEDFAA8EBAC048D2067E5B0158325F
(sCD3268FB2E69A058B357988C1BAD31C26B18C0D3 - s2B661762AEA08905D55D9C993A5A3B37FF2EC6CD -1 downto 0);  sCBB4558CFEFE324102C5417B1E5A0CBDB858B168(sCD3268FB2E69A058B357988C1BAD31C26B18C0D3 downto sCD3268FB2E69A058B357988C1BAD31C26B18C0D3-8) <= "000000001" ; 
 end if; if s1792FD2BB24BFB0793974D92FA74B345EB0CCAF3 = '1' then  sCBB4558CFEFE324102C5417B1E5A0CBDB858B168 <= '0' & sCBB4558CFEFE324102C5417B1E5A0CBDB858B168 (sCD3268FB2E69A058B357988C1BAD31C26B18C0D3 -2 downto 0) & '0'; end if; if s064596695B62E7458EDC8A508E0EE076015E8499
 = '1' then  sCBB4558CFEFE324102C5417B1E5A0CBDB858B168 <= (others=>'0') ;  if s67A0998548ED967361FBF09931BE2B937104D248 = '1' or s49807CD868D22833D34695DE61B3DA5F68DD41DC = '1' then case sEA8188CAD31707F17B299650F81C67D601FE09D7 is when "001110" | "011100" | "100011" | "101010" | "110001" => 
 sCBB4558CFEFE324102C5417B1E5A0CBDB858B168 (30 downto 0) <= sCBB4558CFEFE324102C5417B1E5A0CBDB858B168 (29 downto 0) & sF4DBC68D16423B9DD337E166EF77471DCEA3D993;  when others =>  sCBB4558CFEFE324102C5417B1E5A0CBDB858B168 <= '0' & sCAF301BC43AEA5B1C0FCEBF9360CAC2EDDDEF3D5
(sCD3268FB2E69A058B357988C1BAD31C26B18C0D3 downto 1);  end case; elsif sCBF7A0249B3E467C859DC6110B4A5C709856666B = '1' or sA8F3D27EFD5141F07A5CE1B87DA29A4ABD9AF24E = '1' then sCBB4558CFEFE324102C5417B1E5A0CBDB858B168 (28 downto 0) <= sCBB4558CFEFE324102C5417B1E5A0CBDB858B168
 (27 downto 0) & sF4DBC68D16423B9DD337E166EF77471DCEA3D993;  elsif sDE7CDC6FDA2463F07579EEEE09153F29DF743435 = '1' or s776F81CD2516996DEA92F16B486A7FED89C09EB8 = '1' then sCBB4558CFEFE324102C5417B1E5A0CBDB858B168 (28 downto 0) <= sCBB4558CFEFE324102C5417B1E5A0CBDB858B168
 (27 downto 0) & sF4DBC68D16423B9DD337E166EF77471DCEA3D993;  end if; if s4045C346006E7236123346044B3C0BBE00D1391F = '1' then  s3C3AD1732E30E3202F031BD11ADED227CB12BDB6 <= sF4DBC68D16423B9DD337E166EF77471DCEA3D993 & s3C3AD1732E30E3202F031BD11ADED227CB12BDB6
 (4 downto 1);  end if; end if; end if; end if; end process; s1792FD2BB24BFB0793974D92FA74B345EB0CCAF3 <= s3DE9704ED5E8C46005ACD085579D848AC14D5B18 and s3878B21E042F1AD8CD97DB6E7D00908A99649D03 and (s0C95BB05F974B637452566ABF145558806623663 or s6A18EECF6FABFF8383A93194D7C565C57343844A
); s2324B84C04CC4C838C23EB219AAB9CF288E9F546 <= s01AF22A3811BAB6264C575A96A22B593A64576AE and not sAA4741C86EC7F1A9388F089FDAFF07D1332CA196 and s134B4B78A794B9AC71D2041279723343FA183008; s064596695B62E7458EDC8A508E0EE076015E8499 <= s2324B84C04CC4C838C23EB219AAB9CF288E9F546
;                              process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, sA871AC5299DD9A2B5922B93C415099F5B17A2CAA, s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9, s7DC4BA5492A3997AE8E131EA0BD60F3CED572BBD) begin if rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F
) then if sF1FC47B36F2DA843714A618883F345968A471A76 = '0' then s46B3B4D75B1901ADCD5C39F1B58D398BB213B6BF <= '0'; else if s7DC4BA5492A3997AE8E131EA0BD60F3CED572BBD = '1' and s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 = CONV_STD_LOGIC_VECTOR(s11183BFF0C2D855AEA5F48EC192129844E5C157D
, sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81) and sA871AC5299DD9A2B5922B93C415099F5B17A2CAA = "0101" then s46B3B4D75B1901ADCD5C39F1B58D398BB213B6BF <= '1'; end if; if s48925532037BE5F8C053A6D5DB7767BB7A703DCF = '1' then s46B3B4D75B1901ADCD5C39F1B58D398BB213B6BF
 <= '0'; end if; end if; end if; end process; s48925532037BE5F8C053A6D5DB7767BB7A703DCF <= '1' when s01AF22A3811BAB6264C575A96A22B593A64576AE = '1' and sAA4741C86EC7F1A9388F089FDAFF07D1332CA196 = '0' and s46B3B4D75B1901ADCD5C39F1B58D398BB213B6BF = '1' else
 '0';  process(s82C78E3CD667612DE97ED7C5FA8365F21045093F) begin if rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then if sF1FC47B36F2DA843714A618883F345968A471A76 = '0' then s035B34BD1D4E71D6E05E7E0C12748A22F2AB0BAF <= '0'; s134B4B78A794B9AC71D2041279723343FA183008
 <= '0'; else s035B34BD1D4E71D6E05E7E0C12748A22F2AB0BAF <= s134B4B78A794B9AC71D2041279723343FA183008; if sA871AC5299DD9A2B5922B93C415099F5B17A2CAA = "0101" then if s48925532037BE5F8C053A6D5DB7767BB7A703DCF = '1' then s134B4B78A794B9AC71D2041279723343FA183008
 <= '1'; end if; elsif sA871AC5299DD9A2B5922B93C415099F5B17A2CAA = "1111" or sA871AC5299DD9A2B5922B93C415099F5B17A2CAA = "1010" then s134B4B78A794B9AC71D2041279723343FA183008 <= '0'; end if; end if; end if; end process;                     s8507177FCFDBD094828F65353CFC1170B6FEA614
 <= s2324B84C04CC4C838C23EB219AAB9CF288E9F546 and sC1AA6E43EDA79EA468391A422C8C0A84CAFE4DD9; sD3C21919EB55E97996C06C9C04A4B4F55DB44A0B <= s8507177FCFDBD094828F65353CFC1170B6FEA614; s27D6EF4CA3309F1B892E6207A8D14DCC6F949466 <= '0' when s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9
 = CONV_STD_LOGIC_VECTOR(s11183BFF0C2D855AEA5F48EC192129844E5C157D, sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81) else  '0' when s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 < CONV_STD_LOGIC_VECTOR( 5, sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81) else (s67A0998548ED967361FBF09931BE2B937104D248
 and s134B4B78A794B9AC71D2041279723343FA183008); s4045C346006E7236123346044B3C0BBE00D1391F <= '1' when (s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 < CONV_STD_LOGIC_VECTOR( 5, sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81)) else '0';  s63DCD945122E83C803DEB91867786995FFCFE62A
 <= '0' when s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 = CONV_STD_LOGIC_VECTOR(29, sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81) else  '0' when s4E7BDE5B3AB15C13905C9F70B630AE314A1BD6A9 < CONV_STD_LOGIC_VECTOR( 5, sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81) else
 ((sCBF7A0249B3E467C859DC6110B4A5C709856666B or sDE7CDC6FDA2463F07579EEEE09153F29DF743435) and s134B4B78A794B9AC71D2041279723343FA183008); sC1AA6E43EDA79EA468391A422C8C0A84CAFE4DD9 <= s63DCD945122E83C803DEB91867786995FFCFE62A when sA871AC5299DD9A2B5922B93C415099F5B17A2CAA
 = "1000" else  s63DCD945122E83C803DEB91867786995FFCFE62A when sA871AC5299DD9A2B5922B93C415099F5B17A2CAA = "1001" else  s27D6EF4CA3309F1B892E6207A8D14DCC6F949466; s78D1CF9FDB871B9B4256DCE09B67D406079A5FB8 <= ((sD3C21919EB55E97996C06C9C04A4B4F55DB44A0B and
 s9606968BB22D6E6CABE7FC03219FFECDA4CB919D(4)) xor sF4DBC68D16423B9DD337E166EF77471DCEA3D993); process(s82C78E3CD667612DE97ED7C5FA8365F21045093F) begin if rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then if (sF1FC47B36F2DA843714A618883F345968A471A76
 = '0') then s9606968BB22D6E6CABE7FC03219FFECDA4CB919D <= "11111"; else if s86F6EB29E2D65A736372F43D1F449BCF6DB2BA0A ='1' or s34D0BA0417C5C46CBC3249708B1E4BB573BE4F13 ='1' or s3B95BCD02DFA6D86D669FA75993367A9B3D3207A ='1' then s9606968BB22D6E6CABE7FC03219FFECDA4CB919D
 <= "11111"; elsif (sD3C21919EB55E97996C06C9C04A4B4F55DB44A0B ='1') then s9606968BB22D6E6CABE7FC03219FFECDA4CB919D(4) <= s9606968BB22D6E6CABE7FC03219FFECDA4CB919D(3); s9606968BB22D6E6CABE7FC03219FFECDA4CB919D(3) <= ((s78D1CF9FDB871B9B4256DCE09B67D406079A5FB8
 and sD3C21919EB55E97996C06C9C04A4B4F55DB44A0B) xor s9606968BB22D6E6CABE7FC03219FFECDA4CB919D(2)); s9606968BB22D6E6CABE7FC03219FFECDA4CB919D(2) <= s9606968BB22D6E6CABE7FC03219FFECDA4CB919D(1); s9606968BB22D6E6CABE7FC03219FFECDA4CB919D(1) <= ((s78D1CF9FDB871B9B4256DCE09B67D406079A5FB8
 and sD3C21919EB55E97996C06C9C04A4B4F55DB44A0B) xor s9606968BB22D6E6CABE7FC03219FFECDA4CB919D(0)); s9606968BB22D6E6CABE7FC03219FFECDA4CB919D(0) <= s78D1CF9FDB871B9B4256DCE09B67D406079A5FB8; end if; end if; end if; end process; s0BFFA2AEF006C5821760F1A640F5456669E1486A
 <= '1' when ((s74009442A8C13802B71EA10AB67B2A147A944F36 /= s228AB3A49C983930DA44D78299DB703391BE79F3) and (s34D0BA0417C5C46CBC3249708B1E4BB573BE4F13 = '1' or s3B95BCD02DFA6D86D669FA75993367A9B3D3207A = '1' or s855750D5D93589BB5ABD95DCDECD97BED3D7389E = '1')) else '0'; s74009442A8C13802B71EA10AB67B2A147A944F36 <= s3C3AD1732E30E3202F031BD11ADED227CB12BDB6(0) & s3C3AD1732E30E3202F031BD11ADED227CB12BDB6(1) & s3C3AD1732E30E3202F031BD11ADED227CB12BDB6(2) & s3C3AD1732E30E3202F031BD11ADED227CB12BDB6(3) & s3C3AD1732E30E3202F031BD11ADED227CB12BDB6
(4); s43F7D19F6FFB52EF969FC2858BC1CA57C001562A <= s74009442A8C13802B71EA10AB67B2A147A944F36; s228AB3A49C983930DA44D78299DB703391BE79F3 <= not s9606968BB22D6E6CABE7FC03219FFECDA4CB919D(4 downto 0); sEA8188CAD31707F17B299650F81C67D601FE09D7 <= sE420A02AD972A785E332BF27D04B53B8868A4F0E
 (29 downto 24);  process(s82C78E3CD667612DE97ED7C5FA8365F21045093F) begin if rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then if sF1FC47B36F2DA843714A618883F345968A471A76 = '0' then s013E9FFBF04A31B71784E98EAB7A683996BA039E <= (others => '0'); sBE3694D6DE3020DED7EF579482C5628CB0A7D85D <= '0'; s9279E19351BBF8CD9801F2005A998BF5C72988B9 <= '0'; s34D0BA0417C5C46CBC3249708B1E4BB573BE4F13 <= '0'; s3B95BCD02DFA6D86D669FA75993367A9B3D3207A <= '0'; s855750D5D93589BB5ABD95DCDECD97BED3D7389E <= '0'; s298D55696DC353303493AAE18ABFD0C95B97F0F7
 <= '1'; else s34D0BA0417C5C46CBC3249708B1E4BB573BE4F13 <= s03384791D53DA7C796CA8B60E2BF84B83EF294E1; s3B95BCD02DFA6D86D669FA75993367A9B3D3207A <= s3FE6E74D86F2DF0268B67C717D22E60D521CE7E5; s855750D5D93589BB5ABD95DCDECD97BED3D7389E <= sD02015CB26E1B7025DF2F7880CFEB9376D504E69
; s298D55696DC353303493AAE18ABFD0C95B97F0F7 <= s8949CFA6A16FC99FBD129BE88F26A12A41A2ACE1; case sEA8188CAD31707F17B299650F81C67D601FE09D7 is when "000111" =>  if s03384791D53DA7C796CA8B60E2BF84B83EF294E1 = '1' then s013E9FFBF04A31B71784E98EAB7A683996BA039E
 <= ('0' & sCBB4558CFEFE324102C5417B1E5A0CBDB858B168(sCD3268FB2E69A058B357988C1BAD31C26B18C0D3 -1 downto 1)); sBE3694D6DE3020DED7EF579482C5628CB0A7D85D <= sCBB4558CFEFE324102C5417B1E5A0CBDB858B168(0); s9279E19351BBF8CD9801F2005A998BF5C72988B9 <= '0'; end 
if; when "111000" | "001001" | "011011" | "100100" | "101101" | "110110" =>  if s03384791D53DA7C796CA8B60E2BF84B83EF294E1 = '1' then s013E9FFBF04A31B71784E98EAB7A683996BA039E <= ("00" & sCBB4558CFEFE324102C5417B1E5A0CBDB858B168(sCD3268FB2E69A058B357988C1BAD31C26B18C0D3
 -1 downto 2)); sBE3694D6DE3020DED7EF579482C5628CB0A7D85D <= sCBB4558CFEFE324102C5417B1E5A0CBDB858B168(0); s9279E19351BBF8CD9801F2005A998BF5C72988B9 <= not sCBB4558CFEFE324102C5417B1E5A0CBDB858B168(1); end if; when others =>  if s03384791D53DA7C796CA8B60E2BF84B83EF294E1
 = '1' then s013E9FFBF04A31B71784E98EAB7A683996BA039E <= ("00000" & sCBB4558CFEFE324102C5417B1E5A0CBDB858B168(sCD3268FB2E69A058B357988C1BAD31C26B18C0D3 -1 downto 5)); sBE3694D6DE3020DED7EF579482C5628CB0A7D85D <= '0'; s9279E19351BBF8CD9801F2005A998BF5C72988B9
 <= '0'; end if; end case; if s3FE6E74D86F2DF0268B67C717D22E60D521CE7E5 = '1' or sD02015CB26E1B7025DF2F7880CFEB9376D504E69 = '1' then  s013E9FFBF04A31B71784E98EAB7A683996BA039E <= ("00000" & sCBB4558CFEFE324102C5417B1E5A0CBDB858B168(sCD3268FB2E69A058B357988C1BAD31C26B18C0D3
 -1 downto 5)); end if; end if; end if; end process;  process(sEA8188CAD31707F17B299650F81C67D601FE09D7) begin case sEA8188CAD31707F17B299650F81C67D601FE09D7 is when "001001" | "011011" | "100100" | "101101" | "110110" =>  sA73098C7B13AE4EE2D18DD1A3C28A605F0315F7B
 <= '1'; when others => sA73098C7B13AE4EE2D18DD1A3C28A605F0315F7B <= '0'; end case; end process; s8949CFA6A16FC99FBD129BE88F26A12A41A2ACE1 <= '0' when sA73098C7B13AE4EE2D18DD1A3C28A605F0315F7B = '1' and sA871AC5299DD9A2B5922B93C415099F5B17A2CAA = "0101" and
 sC95BB2A3A95288115289D986565E400E04F2B5A0 = '1' else  '0' when sA73098C7B13AE4EE2D18DD1A3C28A605F0315F7B = '1' and sA871AC5299DD9A2B5922B93C415099F5B17A2CAA = "1000" and sC95BB2A3A95288115289D986565E400E04F2B5A0 = '1' else  '0' when sA73098C7B13AE4EE2D18DD1A3C28A605F0315F7B
 = '1' and sA871AC5299DD9A2B5922B93C415099F5B17A2CAA = "1001" and sC95BB2A3A95288115289D986565E400E04F2B5A0 = '1' else  '0' when sA73098C7B13AE4EE2D18DD1A3C28A605F0315F7B = '1' and sA871AC5299DD9A2B5922B93C415099F5B17A2CAA = "1010" and sC95BB2A3A95288115289D986565E400E04F2B5A0
 = '1' else  '0' when sA73098C7B13AE4EE2D18DD1A3C28A605F0315F7B = '1' and sA871AC5299DD9A2B5922B93C415099F5B17A2CAA = "1011" and sC95BB2A3A95288115289D986565E400E04F2B5A0 = '1' else  s3878B21E042F1AD8CD97DB6E7D00908A99649D03 when sA73098C7B13AE4EE2D18DD1A3C28A605F0315F7B
 = '1' and sA871AC5299DD9A2B5922B93C415099F5B17A2CAA > "1011" else  s73124B1BDDFA8E0A4B7A0970B215A0C89FD997AA; s1504ADD95BA0488B2CA487398BBC3A3FB56ED3A4 <= sD24BF1A9310E03CA3B5DBECC807B894C04E87F42; s858AFDE712A6913772203E81B3BDEEB1165DDD96 <= sCBB4558CFEFE324102C5417B1E5A0CBDB858B168
(sCD3268FB2E69A058B357988C1BAD31C26B18C0D3 -5) when sA73098C7B13AE4EE2D18DD1A3C28A605F0315F7B = '1' and sA871AC5299DD9A2B5922B93C415099F5B17A2CAA > "1001" else  sCBB4558CFEFE324102C5417B1E5A0CBDB858B168(sCD3268FB2E69A058B357988C1BAD31C26B18C0D3 -1) when sA871AC5299DD9A2B5922B93C415099F5B17A2CAA
 = "0001" else '0'; s1FAAEBEE7B845D3CBACD553CA078AD4D43E0ADFA <= s035B34BD1D4E71D6E05E7E0C12748A22F2AB0BAF and (not s134B4B78A794B9AC71D2041279723343FA183008); s03384791D53DA7C796CA8B60E2BF84B83EF294E1 <= (sA8F3D27EFD5141F07A5CE1B87DA29A4ABD9AF24E and (not
 s69B82088412476FAF1B1D1362493AAF169716766 )) when s90196555A8BFC1A5EE5D4925FBA2AF598F9D76F9 = "01" else (sA8F3D27EFD5141F07A5CE1B87DA29A4ABD9AF24E and (not s69B82088412476FAF1B1D1362493AAF169716766 )) when s90196555A8BFC1A5EE5D4925FBA2AF598F9D76F9 = "10" 
else (s1D698942AE29B843C12FC388FE7AE002990CA8DC and (not s7B2460199CAF56FF7F3235463ED56BE379DEF304)) when (s90196555A8BFC1A5EE5D4925FBA2AF598F9D76F9 = "00" and sA73098C7B13AE4EE2D18DD1A3C28A605F0315F7B = '1') else s1FAAEBEE7B845D3CBACD553CA078AD4D43E0ADFA
; s3FE6E74D86F2DF0268B67C717D22E60D521CE7E5 <= (s776F81CD2516996DEA92F16B486A7FED89C09EB8 and (not sA03ED9A8ADD1D6369CFFD09A3B204681F4FD4323)) when s90196555A8BFC1A5EE5D4925FBA2AF598F9D76F9 = "10" else s1FAAEBEE7B845D3CBACD553CA078AD4D43E0ADFA when s90196555A8BFC1A5EE5D4925FBA2AF598F9D76F9
 = "01" else '0'; sD02015CB26E1B7025DF2F7880CFEB9376D504E69 <= s1FAAEBEE7B845D3CBACD553CA078AD4D43E0ADFA when s90196555A8BFC1A5EE5D4925FBA2AF598F9D76F9 = "10" else '0'; s353B8D288425991916C61A5A9DFE44B11BBCF753 <= s013E9FFBF04A31B71784E98EAB7A683996BA039E
; sA16C86782D377069727114AB99F123218DC1EE4E <= s34D0BA0417C5C46CBC3249708B1E4BB573BE4F13; s07A72EEC7FE78460042B89F4D0DA7BE551FEC90A <= s3B95BCD02DFA6D86D669FA75993367A9B3D3207A; s28EDCB4BE5AFFD576E337FA1A3A5AAEEA7D7B33C <= s855750D5D93589BB5ABD95DCDECD97BED3D7389E
; sC4B6EA407C3AA8DD2E6A18E7F77C14FACC951414 <= sBE3694D6DE3020DED7EF579482C5628CB0A7D85D and s34D0BA0417C5C46CBC3249708B1E4BB573BE4F13; s06E676C0BDF7C68FD7495790A14A2FEBA13D3DB6 <= s9279E19351BBF8CD9801F2005A998BF5C72988B9 and s34D0BA0417C5C46CBC3249708B1E4BB573BE4F13
; s32CF03224D0C548C4F44A5420AF0E47F9CE9CB0F <= '1' when s34D0BA0417C5C46CBC3249708B1E4BB573BE4F13 = '1' and (s013E9FFBF04A31B71784E98EAB7A683996BA039E(23 downto 0) = "111111111111111111111111" ) and (s74009442A8C13802B71EA10AB67B2A147A944F36 = "11111") and
 (sEA8188CAD31707F17B299650F81C67D601FE09D7 = "001110" or  sEA8188CAD31707F17B299650F81C67D601FE09D7 = "011100" or  sEA8188CAD31707F17B299650F81C67D601FE09D7 = "100011" or  sEA8188CAD31707F17B299650F81C67D601FE09D7 = "101010" or  sEA8188CAD31707F17B299650F81C67D601FE09D7
 = "110001" or  sEA8188CAD31707F17B299650F81C67D601FE09D7 = "010010")  else '0'; s601E9D380BAA3E6CC5A2AEE58C2C073DF7C885D1 <= '1' when s34D0BA0417C5C46CBC3249708B1E4BB573BE4F13 = '1' and (and_reduce (s013E9FFBF04A31B71784E98EAB7A683996BA039E(23 downto 0) 
xor sE420A02AD972A785E332BF27D04B53B8868A4F0E(23 downto 0)) ='1') and (sEA8188CAD31707F17B299650F81C67D601FE09D7 = "001110" or  sEA8188CAD31707F17B299650F81C67D601FE09D7 = "011100" or  sEA8188CAD31707F17B299650F81C67D601FE09D7 = "100011" or  sEA8188CAD31707F17B299650F81C67D601FE09D7
 = "101010" or  sEA8188CAD31707F17B299650F81C67D601FE09D7 = "110001" or  sEA8188CAD31707F17B299650F81C67D601FE09D7 = "010010")  else '0'; sA516DA7C751934DBE51FECC222FA4984B32B3692 <= '1' when s3B95BCD02DFA6D86D669FA75993367A9B3D3207A ='1' and s90196555A8BFC1A5EE5D4925FBA2AF598F9D76F9
 = "01" and (s013E9FFBF04A31B71784E98EAB7A683996BA039E(20 downto 16) = "01111") else  '1' when s855750D5D93589BB5ABD95DCDECD97BED3D7389E ='1' and s90196555A8BFC1A5EE5D4925FBA2AF598F9D76F9 = "10" and (s013E9FFBF04A31B71784E98EAB7A683996BA039E(20 downto 16) = "01111") 
else  '0'; s7975BCABF4261F33B14B8E6E764BC7741562D89E <= '1' when s3B95BCD02DFA6D86D669FA75993367A9B3D3207A ='1' and s90196555A8BFC1A5EE5D4925FBA2AF598F9D76F9 = "01" and (s013E9FFBF04A31B71784E98EAB7A683996BA039E(20 downto 16) = "11111") else  '1' when s3B95BCD02DFA6D86D669FA75993367A9B3D3207A
 ='1' and s90196555A8BFC1A5EE5D4925FBA2AF598F9D76F9 = "10" and (s013E9FFBF04A31B71784E98EAB7A683996BA039E(20 downto 16) = "11111") else  '0'; s8ABB29C3748C74A80027187254C15F46F51EF2A2 <= sA871AC5299DD9A2B5922B93C415099F5B17A2CAA; s83F675DB784B205945DE32DEA0270B2CF41801FE
 <= s3943BBC49DABABC540DBFCA8F53E255877F4D8F1;  sEE9824B19D5949D38E7E218C1709BFC0B6FFDF6E : pdm generic map( s8012194BD35F0878CACF167A77EE7A04F42ED698 => 10,  s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95 => s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95,   s4A8616F7DBB06E84D521DFE24490E8ADB037CBB1
 => s4A8616F7DBB06E84D521DFE24490E8ADB037CBB1,  s745F184CD6754435326632E8F885833C3FD28CAA => s745F184CD6754435326632E8F885833C3FD28CAA)  port map ( s82C78E3CD667612DE97ED7C5FA8365F21045093F => s82C78E3CD667612DE97ED7C5FA8365F21045093F,  sF1FC47B36F2DA843714A618883F345968A471A76
 => sF1FC47B36F2DA843714A618883F345968A471A76,   sA73098C7B13AE4EE2D18DD1A3C28A605F0315F7B => sA73098C7B13AE4EE2D18DD1A3C28A605F0315F7B,  s90196555A8BFC1A5EE5D4925FBA2AF598F9D76F9 => s90196555A8BFC1A5EE5D4925FBA2AF598F9D76F9,  pdm => s6A5FE1CD0E944495E6BF7242D05EAEACFBA89ACF
,  sA871AC5299DD9A2B5922B93C415099F5B17A2CAA => sA871AC5299DD9A2B5922B93C415099F5B17A2CAA,  s3DE9704ED5E8C46005ACD085579D848AC14D5B18 => s3DE9704ED5E8C46005ACD085579D848AC14D5B18,  s3878B21E042F1AD8CD97DB6E7D00908A99649D03 => s3878B21E042F1AD8CD97DB6E7D00908A99649D03
,  s134B4B78A794B9AC71D2041279723343FA183008 => s134B4B78A794B9AC71D2041279723343FA183008,  s264475A303AC7031FBC8591205A50743DAEAD9CA => sF4DBC68D16423B9DD337E166EF77471DCEA3D993,  s125623D1F098599393E5DE6A762EFFC9DACED467 => s125623D1F098599393E5DE6A762EFFC9DACED467
,  s3943BBC49DABABC540DBFCA8F53E255877F4D8F1 => s3943BBC49DABABC540DBFCA8F53E255877F4D8F1,  sC95BB2A3A95288115289D986565E400E04F2B5A0 => sC95BB2A3A95288115289D986565E400E04F2B5A0,  s79CBDE1F1AE76DE1CEAD5B67EFDA2C6953987F5C => sAA4741C86EC7F1A9388F089FDAFF07D1332CA196
,  sEA5E54196582D991021F5AB19DAC58C70947FB22 => sE734111027AE4A3C909A98A63E7589D18CBEA161, s1B88525B5C44F4D86E63397D61F66E7B1225355E => s1B88525B5C44F4D86E63397D61F66E7B1225355E,   s11183BFF0C2D855AEA5F48EC192129844E5C157D => s11183BFF0C2D855AEA5F48EC192129844E5C157D
 ,  s940FAE140F86D7AAE5446A4FA8C953A8EA6B637D => s0572647003D0AE885FEB3E9760C0F5C78BA6B52A  );  end s75BE5DEF24CA4A61B9676CCF1CC90EBA505DC89E;          