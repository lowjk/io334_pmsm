library ieee; use ieee.std_logic_1164.all; use ieee.numeric_std.all; entity BISS_control is port ( s82C78E3CD667612DE97ED7C5FA8365F21045093F : in std_logic; s0A61EC3B284D41A7527B973B71395AF396BD0749 : in std_logic; sEC9D498A27032D5D5CC9FBE9786A936DA84A5766
 : in std_logic; sADBC8E7E04FA85F5322F3AAA6BF0398152DF9E93 : in std_logic; s67AA1F47031AD081937F209C8CEB3917E3285B98 : in std_logic; sBF63B84FE256F013F6F36AB8B222082B8647B811 : in std_logic_vector(7 downto 0);  s865C7DE113F62D5D7CAC52C2E96B9519EB8FF306 : 
in std_logic_vector(15 downto 0); sE9D5A330018FD42F21BED92AE3F25BEBD3119C81 : out std_logic; s8D52A510B7F21BBB60B0674B11C3DA67D5DE5713 : out std_logic; s6C6651D383B41FAFDF50F2BAA251FDC2A08AB191 : out std_logic; s4F8467F3FA446F57411E855E04FB8C5F7C144A28 : 
out std_logic_vector(63 downto 0); sE4ED7921C578950CCEB828999E51D6DAE12F5A90 : out std_logic;  s4088069AAB16D293A7469FD360A0287D49DE79AE : in std_logic; s76D10F4B556F2B64C06E85300CE7EC78B730048A : in std_logic ); end BISS_control; architecture rtl of BISS_control
 is  type sA564510C7FCE7940D7D16C6D98FB4EC28EF9532B is (s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C, s42904902893D86F1F96274B293D894D00B90EC0C, sA5404BDB4E3CB8663F97DD6FB83BA2227495D22D, sAA38BDF3533DD3CDECA8AAE2000D63F786654426, sCDBEF1C39E592D9A3DD3AD96ED3E14C04C71089A
, sE02D13964AAA0AFC4D9B66B8F5F927AAACD04179, s5FEBF388F22BCBEA400B11D565AA40015BAA27BA, sA8C162BE66CA9216071F4DD4FE349F9E01B4C392, s7A1CA9723971E9E09C282CBEF5151C2B94D35A6C, s22C8A9EFA393E2CC132E38563AE1D741D059113D, s0EE8FCB0FDF901D9B0D26793C62DE7FCC0085E3D
, sFB5597E6B426CF55EEE53274AC5891E98DBCEE79, sE0E4F2883171C2D3103F9C5E105BE2796C1D0D20, s9AEE4C17C38159EB8E63E2146A2FBF6255DB53A4, s9F74852C360D0731C4A69BB7F9C9B6180BA9AFEE); signal sF1D6856D8C6E7F12EED89D6F5F90C7580EF3FE5E, sC3F360CDD6D534EE7E5EB80085F8A784CFE01687
 : sA564510C7FCE7940D7D16C6D98FB4EC28EF9532B;  signal s4729D72C983E68611F3D2F170962E438D6EEC729 : unsigned(15 downto 0); signal s078316AFF6BEB1FA1A2A97CE17D622DE2C01F0AB, sCE4A9CD62E6A2AB3957E4B3743B0900B7E398765 : std_logic;  signal sE8ED6835D5D9F9DB6B1E613C6659B9CB49707489
 : unsigned(9 downto 0); signal s7D421768169CE02634C5F9A247D21A30EB3BA348 : unsigned(15 downto 0); signal s1933CD31C2CAD7E35ECCFB532696A7E6679201C7 : unsigned(7 downto 0); signal s5671B60ACA79D7E7AAA362220DBBEB27307BB408, sF33115B7AD1B39A9F286BD8E6AC7C2B03D8C6771
 : std_logic; signal s5087A156F97E44C8B4FA4E4028F2BE8C50DAA8BD : std_logic; signal s00506246AD19C23077849FB3ED52A1D57EAB8122 : std_logic; signal sE36A0558667B7BAC11863457B94185BFF46FDB4D : std_logic; signal s5724103C905B1DD81E89674E48BBD9329E45720F : std_logic
; signal sFB3107C8B48BCEDD631D98C6FE24FDE2FE5B35FC : std_logic; signal s2EB269661807F704AC7FCE80F96D450960E95BB2, sA63D3E6DF73AB346E87FC63C01AED1D97F96D91D, sD8B326FE5C2DC0FAB305A3EC3CAB5B7338123439 : std_logic; signal s74EEE1FFEA07E4C7E6716BF94B0F961C05D26C62
 : std_logic_vector(2 downto 0); signal sF3E0BFA8E9F591147156A251FCF8ECD8A55B9DEA : std_logic; signal sABECA4F299B2C6E8A00F28EA6D6F8753B3CECD1E : std_logic_vector(1023 downto 0); signal s8DC239BAE0C4B59356AE3036500FFCCDBBFA8E72 : std_logic_vector(63 downto
 0); signal s3D2B651BC6F8DAD148B1D96E9BB80F63FED28E1F, sFD3787837EA190C4D1C4FF997E6A3CBF927B3EDD : std_logic; signal s3CEE9E0D841A89946A317BDFEEDF99D8F9ED8DC0, sF3F5D68E172988078B9E123657D3937649BDABE6 : std_logic; signal s711E1DFE909B9691C0BE2BDD557C4E4D3BE7F06E
, s2CC9648F3BE766AD963F4674275246BB5BDC578E, sB5D8CF0FAC4652151001D86FB268CC6BD905FE47 : std_logic; begin sA0E3F628288F9FF5ED44D93BDADE0807C5D95734 : process(sF1D6856D8C6E7F12EED89D6F5F90C7580EF3FE5E, s67AA1F47031AD081937F209C8CEB3917E3285B98, sF3E0BFA8E9F591147156A251FCF8ECD8A55B9DEA
, sFD3787837EA190C4D1C4FF997E6A3CBF927B3EDD, s3D2B651BC6F8DAD148B1D96E9BB80F63FED28E1F, sADBC8E7E04FA85F5322F3AAA6BF0398152DF9E93, sEC9D498A27032D5D5CC9FBE9786A936DA84A5766, s4729D72C983E68611F3D2F170962E438D6EEC729, sF3F5D68E172988078B9E123657D3937649BDABE6
, s3CEE9E0D841A89946A317BDFEEDF99D8F9ED8DC0, s1933CD31C2CAD7E35ECCFB532696A7E6679201C7, sBF63B84FE256F013F6F36AB8B222082B8647B811, s5087A156F97E44C8B4FA4E4028F2BE8C50DAA8BD) begin  sCE4A9CD62E6A2AB3957E4B3743B0900B7E398765 <= '0'; s078316AFF6BEB1FA1A2A97CE17D622DE2C01F0AB
 <= '0'; sF33115B7AD1B39A9F286BD8E6AC7C2B03D8C6771 <= '0'; s5671B60ACA79D7E7AAA362220DBBEB27307BB408 <= '0'; s00506246AD19C23077849FB3ED52A1D57EAB8122 <= '0'; sE36A0558667B7BAC11863457B94185BFF46FDB4D <= '0'; sE9D5A330018FD42F21BED92AE3F25BEBD3119C81 <= '0'; s8D52A510B7F21BBB60B0674B11C3DA67D5DE5713 <= '0'; s5724103C905B1DD81E89674E48BBD9329E45720F <= '0'; sFB3107C8B48BCEDD631D98C6FE24FDE2FE5B35FC <= '0'; s2EB269661807F704AC7FCE80F96D450960E95BB2 <= '0'; sA63D3E6DF73AB346E87FC63C01AED1D97F96D91D <= '0'; case
 sF1D6856D8C6E7F12EED89D6F5F90C7580EF3FE5E is when s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C => sE36A0558667B7BAC11863457B94185BFF46FDB4D <= '1'; s078316AFF6BEB1FA1A2A97CE17D622DE2C01F0AB <= '1'; s5671B60ACA79D7E7AAA362220DBBEB27307BB408 <= '1'; sFB3107C8B48BCEDD631D98C6FE24FDE2FE5B35FC
 <= '1'; s2EB269661807F704AC7FCE80F96D450960E95BB2 <= '1'; if s67AA1F47031AD081937F209C8CEB3917E3285B98 = '1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s42904902893D86F1F96274B293D894D00B90EC0C; else sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C
; end if; when s42904902893D86F1F96274B293D894D00B90EC0C => sE9D5A330018FD42F21BED92AE3F25BEBD3119C81 <= '1'; if sADBC8E7E04FA85F5322F3AAA6BF0398152DF9E93 = '1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= sA5404BDB4E3CB8663F97DD6FB83BA2227495D22D; else
 sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s42904902893D86F1F96274B293D894D00B90EC0C; end if; when sA5404BDB4E3CB8663F97DD6FB83BA2227495D22D => sCE4A9CD62E6A2AB3957E4B3743B0900B7E398765 <= '1'; if sF3E0BFA8E9F591147156A251FCF8ECD8A55B9DEA = '0' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687
 <= s9F74852C360D0731C4A69BB7F9C9B6180BA9AFEE; elsif s4729D72C983E68611F3D2F170962E438D6EEC729 > 1 then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= sAA38BDF3533DD3CDECA8AAE2000D63F786654426; else sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= sA5404BDB4E3CB8663F97DD6FB83BA2227495D22D
; end if; when sAA38BDF3533DD3CDECA8AAE2000D63F786654426 => sF33115B7AD1B39A9F286BD8E6AC7C2B03D8C6771 <= '1'; if sFD3787837EA190C4D1C4FF997E6A3CBF927B3EDD='1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= sCDBEF1C39E592D9A3DD3AD96ED3E14C04C71089A; elsif
 s5087A156F97E44C8B4FA4E4028F2BE8C50DAA8BD='1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s9F74852C360D0731C4A69BB7F9C9B6180BA9AFEE; else sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= sAA38BDF3533DD3CDECA8AAE2000D63F786654426; end if; when sCDBEF1C39E592D9A3DD3AD96ED3E14C04C71089A
 => if s3D2B651BC6F8DAD148B1D96E9BB80F63FED28E1F='1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= sE02D13964AAA0AFC4D9B66B8F5F927AAACD04179; elsif s5087A156F97E44C8B4FA4E4028F2BE8C50DAA8BD='1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s9F74852C360D0731C4A69BB7F9C9B6180BA9AFEE
; else sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= sCDBEF1C39E592D9A3DD3AD96ED3E14C04C71089A; end if; when sE02D13964AAA0AFC4D9B66B8F5F927AAACD04179 => if sF3F5D68E172988078B9E123657D3937649BDABE6='1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= sA8C162BE66CA9216071F4DD4FE349F9E01B4C392
; else sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= sE02D13964AAA0AFC4D9B66B8F5F927AAACD04179; end if; when sA8C162BE66CA9216071F4DD4FE349F9E01B4C392 => if sF3F5D68E172988078B9E123657D3937649BDABE6='1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s5FEBF388F22BCBEA400B11D565AA40015BAA27BA
; else sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= sA8C162BE66CA9216071F4DD4FE349F9E01B4C392; end if; when s5FEBF388F22BCBEA400B11D565AA40015BAA27BA => if sF3F5D68E172988078B9E123657D3937649BDABE6='1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s7A1CA9723971E9E09C282CBEF5151C2B94D35A6C
; else sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s5FEBF388F22BCBEA400B11D565AA40015BAA27BA; end if; when s7A1CA9723971E9E09C282CBEF5151C2B94D35A6C => s00506246AD19C23077849FB3ED52A1D57EAB8122 <= '1'; if s1933CD31C2CAD7E35ECCFB532696A7E6679201C7 < unsigned
(sBF63B84FE256F013F6F36AB8B222082B8647B811)-1 then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s5FEBF388F22BCBEA400B11D565AA40015BAA27BA; else sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s22C8A9EFA393E2CC132E38563AE1D741D059113D; end if; when s22C8A9EFA393E2CC132E38563AE1D741D059113D
 => if sEC9D498A27032D5D5CC9FBE9786A936DA84A5766='1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s0EE8FCB0FDF901D9B0D26793C62DE7FCC0085E3D; else sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s22C8A9EFA393E2CC132E38563AE1D741D059113D; end if; when s0EE8FCB0FDF901D9B0D26793C62DE7FCC0085E3D
 => s8D52A510B7F21BBB60B0674B11C3DA67D5DE5713 <= '1'; sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= sFB5597E6B426CF55EEE53274AC5891E98DBCEE79; when sFB5597E6B426CF55EEE53274AC5891E98DBCEE79 => if s5087A156F97E44C8B4FA4E4028F2BE8C50DAA8BD='1' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687
 <= sE0E4F2883171C2D3103F9C5E105BE2796C1D0D20; else sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= sFB5597E6B426CF55EEE53274AC5891E98DBCEE79; end if; when sE0E4F2883171C2D3103F9C5E105BE2796C1D0D20 => s5724103C905B1DD81E89674E48BBD9329E45720F <= '1'; sC3F360CDD6D534EE7E5EB80085F8A784CFE01687
 <= s9AEE4C17C38159EB8E63E2146A2FBF6255DB53A4; when s9AEE4C17C38159EB8E63E2146A2FBF6255DB53A4 => if s67AA1F47031AD081937F209C8CEB3917E3285B98='0' then sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C; else sC3F360CDD6D534EE7E5EB80085F8A784CFE01687
 <= s9AEE4C17C38159EB8E63E2146A2FBF6255DB53A4; end if; when s9F74852C360D0731C4A69BB7F9C9B6180BA9AFEE => sA63D3E6DF73AB346E87FC63C01AED1D97F96D91D <= '1'; sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s22C8A9EFA393E2CC132E38563AE1D741D059113D; when others => sC3F360CDD6D534EE7E5EB80085F8A784CFE01687 <= s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C; end case; end process sA0E3F628288F9FF5ED44D93BDADE0807C5D95734;  s01B836CC599AAC170C41C635FD46B72FA2B88119: process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749
) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749 = '1' then sF1D6856D8C6E7F12EED89D6F5F90C7580EF3FE5E <= s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C; elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then sF1D6856D8C6E7F12EED89D6F5F90C7580EF3FE5E
 <= sC3F360CDD6D534EE7E5EB80085F8A784CFE01687; end if; end process s01B836CC599AAC170C41C635FD46B72FA2B88119;  sE108E47002A868BCBC737ABCADAD955D725DF46E: process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749) begin if
 s0A61EC3B284D41A7527B973B71395AF396BD0749 = '1' then s4729D72C983E68611F3D2F170962E438D6EEC729 <= (others => '0'); elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then if s078316AFF6BEB1FA1A2A97CE17D622DE2C01F0AB = '1' then s4729D72C983E68611F3D2F170962E438D6EEC729
 <= (others => '0'); elsif sCE4A9CD62E6A2AB3957E4B3743B0900B7E398765='1' and sEC9D498A27032D5D5CC9FBE9786A936DA84A5766='1' then s4729D72C983E68611F3D2F170962E438D6EEC729 <= s4729D72C983E68611F3D2F170962E438D6EEC729 + 1; end if; end if; end process sE108E47002A868BCBC737ABCADAD955D725DF46E
;  sDE9428F0AC206F4B59BA95C04AAEA3BC2F6ED8F3: process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749 = '1' then sE8ED6835D5D9F9DB6B1E613C6659B9CB49707489 <= (others => '0'); elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then if s5671B60ACA79D7E7AAA362220DBBEB27307BB408 = '1' then sE8ED6835D5D9F9DB6B1E613C6659B9CB49707489 <= (others => '0'); elsif sF33115B7AD1B39A9F286BD8E6AC7C2B03D8C6771='1' and sE8ED6835D5D9F9DB6B1E613C6659B9CB49707489
< "11" & x"FF" then sE8ED6835D5D9F9DB6B1E613C6659B9CB49707489 <= sE8ED6835D5D9F9DB6B1E613C6659B9CB49707489 + 1; end if; end if; end process sDE9428F0AC206F4B59BA95C04AAEA3BC2F6ED8F3;  process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749
) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749 = '1' then s74EEE1FFEA07E4C7E6716BF94B0F961C05D26C62 <= (others => '0'); elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then s74EEE1FFEA07E4C7E6716BF94B0F961C05D26C62 <= s74EEE1FFEA07E4C7E6716BF94B0F961C05D26C62
(1 downto 0) & s76D10F4B556F2B64C06E85300CE7EC78B730048A; end if; end process; sF3E0BFA8E9F591147156A251FCF8ECD8A55B9DEA <= s74EEE1FFEA07E4C7E6716BF94B0F961C05D26C62(2); s3D2B651BC6F8DAD148B1D96E9BB80F63FED28E1F <= '1' when s74EEE1FFEA07E4C7E6716BF94B0F961C05D26C62
(2 downto 1) = "01" else '0'; sFD3787837EA190C4D1C4FF997E6A3CBF927B3EDD <= '1' when s74EEE1FFEA07E4C7E6716BF94B0F961C05D26C62(2 downto 1) = "10" else '0';  process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749) begin
 if s0A61EC3B284D41A7527B973B71395AF396BD0749 = '1' then sABECA4F299B2C6E8A00F28EA6D6F8753B3CECD1E <= (others => '1'); elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then sABECA4F299B2C6E8A00F28EA6D6F8753B3CECD1E <= sABECA4F299B2C6E8A00F28EA6D6F8753B3CECD1E
(1022 downto 0) & s4088069AAB16D293A7469FD360A0287D49DE79AE; end if; end process; sFA2B865AE18456645D99F93763FC2E7BFD7C47B7 : process(sE8ED6835D5D9F9DB6B1E613C6659B9CB49707489, sABECA4F299B2C6E8A00F28EA6D6F8753B3CECD1E) begin for s020F5125771EEEB6F963720A8BB968FCA977AA41
 in 0 to 1023 loop if s020F5125771EEEB6F963720A8BB968FCA977AA41=to_integer(sE8ED6835D5D9F9DB6B1E613C6659B9CB49707489) then s711E1DFE909B9691C0BE2BDD557C4E4D3BE7F06E <= sABECA4F299B2C6E8A00F28EA6D6F8753B3CECD1E(s020F5125771EEEB6F963720A8BB968FCA977AA41); end
 if; end loop; end process sFA2B865AE18456645D99F93763FC2E7BFD7C47B7;  s1DDD5F0829B5CE25CBF9A343410FB0DA516D24D6: process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749
='1' then s2CC9648F3BE766AD963F4674275246BB5BDC578E <= '0'; sB5D8CF0FAC4652151001D86FB268CC6BD905FE47 <= '0'; elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then sB5D8CF0FAC4652151001D86FB268CC6BD905FE47 <= s711E1DFE909B9691C0BE2BDD557C4E4D3BE7F06E
; s2CC9648F3BE766AD963F4674275246BB5BDC578E <= sB5D8CF0FAC4652151001D86FB268CC6BD905FE47; end if; end process s1DDD5F0829B5CE25CBF9A343410FB0DA516D24D6; s3CEE9E0D841A89946A317BDFEEDF99D8F9ED8DC0 <= '1' when s2CC9648F3BE766AD963F4674275246BB5BDC578E='0' and
 sB5D8CF0FAC4652151001D86FB268CC6BD905FE47='1' else '0'; sF3F5D68E172988078B9E123657D3937649BDABE6 <= '1' when s2CC9648F3BE766AD963F4674275246BB5BDC578E='1' and sB5D8CF0FAC4652151001D86FB268CC6BD905FE47='0' else '0';  s5ACBE19798DCEAD883E451C594458D286F102EAD
: process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749 = '1' then s1933CD31C2CAD7E35ECCFB532696A7E6679201C7 <= (others => '0'); elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F
) then if sFB3107C8B48BCEDD631D98C6FE24FDE2FE5B35FC = '1' then s1933CD31C2CAD7E35ECCFB532696A7E6679201C7 <= (others => '0'); elsif s00506246AD19C23077849FB3ED52A1D57EAB8122='1' then s1933CD31C2CAD7E35ECCFB532696A7E6679201C7 <= s1933CD31C2CAD7E35ECCFB532696A7E6679201C7
 + 1; end if; end if; end process s5ACBE19798DCEAD883E451C594458D286F102EAD;  sCC62984C14BE81D9754B7865F8E489AD7AE01782: process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749
 = '1' then s8DC239BAE0C4B59356AE3036500FFCCDBBFA8E72 <= (others => '0'); elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then if sE36A0558667B7BAC11863457B94185BFF46FDB4D = '1' then s8DC239BAE0C4B59356AE3036500FFCCDBBFA8E72 <= (others => '0'); elsif s00506246AD19C23077849FB3ED52A1D57EAB8122='1' then s8DC239BAE0C4B59356AE3036500FFCCDBBFA8E72 <= s8DC239BAE0C4B59356AE3036500FFCCDBBFA8E72(s8DC239BAE0C4B59356AE3036500FFCCDBBFA8E72'left-1 downto 0) & sF3E0BFA8E9F591147156A251FCF8ECD8A55B9DEA; end if
; end if; end process sCC62984C14BE81D9754B7865F8E489AD7AE01782;  s42770BFA3931C7401F0C247E11F10D222438B64C: process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749 = '1' 
then sD8B326FE5C2DC0FAB305A3EC3CAB5B7338123439 <= '0'; elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then if s2EB269661807F704AC7FCE80F96D450960E95BB2 = '1' then sD8B326FE5C2DC0FAB305A3EC3CAB5B7338123439 <= '0'; elsif sA63D3E6DF73AB346E87FC63C01AED1D97F96D91D
='1' then sD8B326FE5C2DC0FAB305A3EC3CAB5B7338123439 <= '1'; end if; end if; end process s42770BFA3931C7401F0C247E11F10D222438B64C;  s40DE9FB8B6E41E9D684E868566180D8E7D566D3F: process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749
) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749 = '1' then sE4ED7921C578950CCEB828999E51D6DAE12F5A90 <= '0'; s4F8467F3FA446F57411E855E04FB8C5F7C144A28 <= (others => '0'); s6C6651D383B41FAFDF50F2BAA251FDC2A08AB191 <= '0'; elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F
) then s6C6651D383B41FAFDF50F2BAA251FDC2A08AB191 <= '0'; if s5724103C905B1DD81E89674E48BBD9329E45720F = '1' then s4F8467F3FA446F57411E855E04FB8C5F7C144A28 <= s8DC239BAE0C4B59356AE3036500FFCCDBBFA8E72; sE4ED7921C578950CCEB828999E51D6DAE12F5A90 <= sD8B326FE5C2DC0FAB305A3EC3CAB5B7338123439
; s6C6651D383B41FAFDF50F2BAA251FDC2A08AB191 <= '1'; end if; end if; end process s40DE9FB8B6E41E9D684E868566180D8E7D566D3F;  sE89B484851192CC4812859B8C19EB7C1BC90F325: process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749
) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749 = '1' then s7D421768169CE02634C5F9A247D21A30EB3BA348 <= (others => '0'); elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then  if sF1D6856D8C6E7F12EED89D6F5F90C7580EF3FE5E /= sC3F360CDD6D534EE7E5EB80085F8A784CFE01687
 then s7D421768169CE02634C5F9A247D21A30EB3BA348 <= (others => '0'); else s7D421768169CE02634C5F9A247D21A30EB3BA348 <= s7D421768169CE02634C5F9A247D21A30EB3BA348 + 1; end if; end if; end process sE89B484851192CC4812859B8C19EB7C1BC90F325; s5087A156F97E44C8B4FA4E4028F2BE8C50DAA8BD
 <= '1' when s7D421768169CE02634C5F9A247D21A30EB3BA348 >= unsigned(s865C7DE113F62D5D7CAC52C2E96B9519EB8FF306) else '0'; end rtl;