library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;
  use work.ENDAT_SNIFFER_pkg.all;

entity ENDAT_SNIFFER is
  port
  (
    clk_i            : in std_logic;
    reset_i          : in std_logic;              
    
    version         : out std_logic_vector(31 downto 0);     
    
    tReset_i         : in std_logic_vector(31 downto 0);  
    numPulPosVal_i   : in std_logic_vector(31 downto 0);  
    distRev_i        : in std_logic_vector(31 downto 0);  
    
    
    dataValid_o      : out std_logic;
    rxPosVal_o       : out std_logic_vector(31 downto 0); 
    numRev_o         : out std_logic_vector(31 downto 0);
    error_o          : out std_logic_vector(31 downto 0);
        
		
    i_serial_clk     : in std_logic;   
    i_serial         : in std_logic    
  );
end ENDAT_SNIFFER;

architecture Struct OF ENDAT_SNIFFER IS constant s31AF80B9B3671B438C161958C96A8305B72EF8B0 : std_logic_vector(55 downto 0) := (others => '0'); constant s93A6A3A936D92717AE7F5510442BDD1FEF22EC32 : std_logic_vector(55 downto 0) := (others => '1'); constant 
sFA993A047EF0E48F00E39634285E74B781D00DBF : unsigned(31 downto 0) := x"00000002"; constant sE5CEEC534B45504250BB0AB9C68F528B4427B4EA : unsigned(31 downto 0) := x"00000006"; constant sF1ACDF194238D93C80C3F56B982846A83ABF8042 : unsigned(31 downto 0) := x"00000008";
 constant s554B052BE2734AB000DFA8E34A6DCD1C5B7F62F3 : unsigned(31 downto 0) := x"00000010";  constant sF18D65E9875B3783D0FD9B8A653B5F0B9BE8AE44 : unsigned(31 downto 0) := x"00000002"; constant s54450457B8FEB0B916F66422DDC28520A6F27D61 : unsigned(31 downto
 0) := x"00000008"; constant s287FEDCA98AA2143D3F527A97C155CE0F210A782 : unsigned(31 downto 0) := x"00000005";  constant s48ABDA14A8459879C068D03E11C2A85FEBF56F62 : std_logic_vector(31 downto 0) := x"00091050";  constant s10694D6404BE82E7D38125D4E95817256BF8F802
 : std_logic_vector(31 downto 0) := x"00010000";  constant s306BFF0CDBF6BF07A6F7DBB40262760A4BE39DB7 : std_logic_vector(31 downto 0) := x"00000008";   signal s7D425144B574080EAE524904A8A3A1B003EE34A7 : unsigned(31 downto 0); signal sA0F87C252F9449120B37FA8565AD3B246A3EBC17
 : unsigned(31 downto 0); signal sF073296EFBB46BD30ADC8EA25E1CC93687EBDAFB : integer range 0 to 56; type s84A58935577AFA37FF091033F9FB65ACBEB81483 is (s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C, sBB12D33790A5D3018B4D986F4ADB83977C5D8601, s36AC7A0A1A83247FFEBA473A089671A1570A444F
, s4D060726C033C2FAEAF8BEA001EE62AE7781F8FF, s4BD5B45FED6CFDC9C7C9EB134B11243E9E183FB8, s3F5CD917DD715D35070C12A524859CBA336A5E8F, s39F04C15DE0E5F43C559F3657FACB1AA3D4A2CF7, sC4E33B939FA9CAB7BA08E4FBF3DEF9689B5FB0C0, sAC14180D3920A14E53EB388154EEB3BD8EE00F38
, sA265FC1FF568154C90487807499F4E4714E828D2, sA8AD75438F0C3D62010B98FEDD21D5B11EF0BBC1, s529B4ABD50A0DC309F792EE5D475A66D0D9959A2, s4E6FE1CA131098FC04443D071866EADE68B517F4); signal s22E923CF436A1BF1EAA149BF66A7AD165ABABD9A, s2A4FD558F206D02C009EE8C6C3270121218EBF72
 : s84A58935577AFA37FF091033F9FB65ACBEB81483; signal s38B47F4C3DE0DCB215428A00C075B72E81724995, s7BA0158498624EFFF7A85F2DE562B881D380F526 : unsigned(31 downto 0); signal s42C156E01C093831B32D6A7CBFD3020F1F90D4CF : std_logic; signal s1A1FBAC4E57E71A08D58F34D3F236E10FDBB13F1
 : std_logic; signal s8DC239BAE0C4B59356AE3036500FFCCDBBFA8E72 : std_logic; signal s299A4649AF76D252E8BCE9B9976634617E034DC3 : unsigned(31 downto 0); signal s0465AAD501BCFB42A3CE710255F7BF6B54E619DD : std_logic_vector(55 downto 0); signal s9216F1816ACE78FB0851459E9601420ABC3AA570
 : std_logic_vector(1 downto 0); signal s4F8EEACE44418C026D8F7B6609F95D9F2983F61C, sEB2C0A31F86ED13FF0CDECB77CA291A86128B247 : std_logic; signal s2C546333D09386C1C9D785047A9CEA69F8B26C94 : std_logic_vector(4 downto 0); signal s743EE1FDAFD422AABFC09E9E393850C4C85EAD2E
 : std_logic;  signal s0FFAB4F8912FCE63B3997867066DFB9C1F628974, s3538966AA1D4ACE62D812FC8AB90B6A47190487F : std_logic; signal s327A67E98B0309EF07AAC0342DBE9324EEC837C9 : std_logic_vector(127 downto 0); signal s45D2033B63004B619AF223745CE9944CA468D689 : std_logic
; signal sEA8188CAD31707F17B299650F81C67D601FE09D7 : std_logic_vector(5 downto 0); signal s2DE53BABF9E8291149A3F55C3450649370E3009F : std_logic_vector(7 downto 0); signal sDF9F3E40D3B907510D4DF16BCDAFC2586EB30618 : std_logic_vector(15 downto 0); signal sEBDD504D1ED5866A72788C09CE264D16E1872EDC
, s57AE96E3A4322EF36A1E1352A866E15B3C188F64 : std_logic; signal s373038E3F2FB6ECFC8FEB465BD78F4377C39923A, sC3ADFA536EF4E4699F020FEC7F3F5E5F95645E71 : std_logic; signal s395EF2527A3109AD4086230A8FD7F23B1F2F0F41 : std_logic; signal s08140CA014D79009968544D9ECD7EAA0E163EED4
 : std_logic; signal s2F285CF0B57A3B502B36C687EFD83233AC8934DC : unsigned(31 downto 0); signal s9E27824C43FC3BC94286CC02E57D7EA018AB2D12 : unsigned(31 downto 0); signal sA2DAE05A577AC12D23A3CED89B449A366DCFF9D3 : unsigned(31 downto 0); signal s1E9AD3357247BE14ACDD8BA1FE752CC280C75D49
 : std_logic; signal s2352BDBE6CE03BBCE38F2DE675BB47F601C0CEE4 : std_logic; signal sDEB77204C753BE668599CE98F2768D24342B4D6B, s44987DF76FE68D9CEF103968757796A160C63E1C : std_logic; signal s803DC9CAA8B495BF1BF7AC678ABDB7265B406E97, s8E9F68EAF8B9CC6752ACCB89FC9C7B7337F6BBA7
 : std_logic; signal s5960FAE099FE1D30E1893ED128A9BC168134F816 : std_logic; constant s18232216D466596BEB636EEAE873919D97A90393 : integer := 32;  signal sB3A8B19CA98570BA8D1B96F098A8058070AA0E06 : integer range 0 to s18232216D466596BEB636EEAE873919D97A90393
;    constant sAD571A7EC29F4958A6460F21AC21EB618B3EAFA0 : integer := 32;  signal s1ECA68304446F3295D7FC3C5B314ADBA0067C044 : integer range 0 to sAD571A7EC29F4958A6460F21AC21EB618B3EAFA0;  signal s38FBA08FA1E8936955F6D21A792256E3658F8387 : std_logic_vector
(31 downto 0);  signal s6D8E140706515F7AFC288159A5BC35A838C23C32 : std_logic_vector(31 downto 0); begin version <= "10" & s731A256AA7EC109FE962BF102445534C5772925D & s7EC4167F3F7F1E99D074313BF18FF4BA05E7ED10 & s5907A17D8E29C7EB61D4F347241BFE4DAC407AEA;  sB3DEBC4A1333AD928E577F918D84173520930691
 : process(clk_i) begin if rising_edge(clk_i) then sEBDD504D1ED5866A72788C09CE264D16E1872EDC <= i_serial_clk; s57AE96E3A4322EF36A1E1352A866E15B3C188F64 <= sEBDD504D1ED5866A72788C09CE264D16E1872EDC; s743EE1FDAFD422AABFC09E9E393850C4C85EAD2E <= s57AE96E3A4322EF36A1E1352A866E15B3C188F64
; end if; end process sB3DEBC4A1333AD928E577F918D84173520930691; s0FFAB4F8912FCE63B3997867066DFB9C1F628974 <= '1' when s743EE1FDAFD422AABFC09E9E393850C4C85EAD2E='0' and s57AE96E3A4322EF36A1E1352A866E15B3C188F64='1' else '0'; s3538966AA1D4ACE62D812FC8AB90B6A47190487F
 <= '1' when s743EE1FDAFD422AABFC09E9E393850C4C85EAD2E='1' and s57AE96E3A4322EF36A1E1352A866E15B3C188F64='0' else '0';  process(clk_i) begin if rising_edge(clk_i) then if reset_i = '1' then s327A67E98B0309EF07AAC0342DBE9324EEC837C9 <= (others => '0'); else
 s327A67E98B0309EF07AAC0342DBE9324EEC837C9 <= s327A67E98B0309EF07AAC0342DBE9324EEC837C9(126 downto 0) & s3538966AA1D4ACE62D812FC8AB90B6A47190487F; end if; end if; end process; s9116D76F37FA5EAA978621D829EEBB6CB2738F91 : process(sA2DAE05A577AC12D23A3CED89B449A366DCFF9D3
, s327A67E98B0309EF07AAC0342DBE9324EEC837C9) begin for s020F5125771EEEB6F963720A8BB968FCA977AA41 in 0 to 127 loop if s020F5125771EEEB6F963720A8BB968FCA977AA41=to_integer(sA2DAE05A577AC12D23A3CED89B449A366DCFF9D3) then s45D2033B63004B619AF223745CE9944CA468D689
 <= s327A67E98B0309EF07AAC0342DBE9324EEC837C9(s020F5125771EEEB6F963720A8BB968FCA977AA41); end if; end loop; end process s9116D76F37FA5EAA978621D829EEBB6CB2738F91;  sDE9E0814E82DB268187B9C25E9114075DCB837C0 : process(clk_i) begin if rising_edge(clk_i) then
 s373038E3F2FB6ECFC8FEB465BD78F4377C39923A <= i_serial; sC3ADFA536EF4E4699F020FEC7F3F5E5F95645E71 <= s373038E3F2FB6ECFC8FEB465BD78F4377C39923A; s395EF2527A3109AD4086230A8FD7F23B1F2F0F41 <= sC3ADFA536EF4E4699F020FEC7F3F5E5F95645E71; end if; end process sDE9E0814E82DB268187B9C25E9114075DCB837C0
;  sA61E52C60F537891176EAE963E0E85484FF304AD : process (clk_i) begin if rising_edge(clk_i) then if reset_i='1' then s22E923CF436A1BF1EAA149BF66A7AD165ABABD9A <= s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C; else s22E923CF436A1BF1EAA149BF66A7AD165ABABD9A <= s2A4FD558F206D02C009EE8C6C3270121218EBF72
; end if; end if; end process sA61E52C60F537891176EAE963E0E85484FF304AD;  s16A54A799612DE170F8EC9B0B99BAC7A233D1DF9 : process(s22E923CF436A1BF1EAA149BF66A7AD165ABABD9A, s2352BDBE6CE03BBCE38F2DE675BB47F601C0CEE4, s395EF2527A3109AD4086230A8FD7F23B1F2F0F41, 
s7BA0158498624EFFF7A85F2DE562B881D380F526, s3538966AA1D4ACE62D812FC8AB90B6A47190487F, s45D2033B63004B619AF223745CE9944CA468D689, s0FFAB4F8912FCE63B3997867066DFB9C1F628974, s42C156E01C093831B32D6A7CBFD3020F1F90D4CF, s38B47F4C3DE0DCB215428A00C075B72E81724995
, s7D425144B574080EAE524904A8A3A1B003EE34A7, s803DC9CAA8B495BF1BF7AC678ABDB7265B406E97, s299A4649AF76D252E8BCE9B9976634617E034DC3) begin  s1A1FBAC4E57E71A08D58F34D3F236E10FDBB13F1 <= '0'; s8DC239BAE0C4B59356AE3036500FFCCDBBFA8E72 <= '0'; case s22E923CF436A1BF1EAA149BF66A7AD165ABABD9A
 is when s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C => if s3538966AA1D4ACE62D812FC8AB90B6A47190487F = '1' then s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= sBB12D33790A5D3018B4D986F4ADB83977C5D8601; else s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C
; end if; when sBB12D33790A5D3018B4D986F4ADB83977C5D8601 => if s38B47F4C3DE0DCB215428A00C075B72E81724995 >= sFA993A047EF0E48F00E39634285E74B781D00DBF then s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s36AC7A0A1A83247FFEBA473A089671A1570A444F; elsif s2352BDBE6CE03BBCE38F2DE675BB47F601C0CEE4
 = '1' then s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s4E6FE1CA131098FC04443D071866EADE68B517F4; else s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= sBB12D33790A5D3018B4D986F4ADB83977C5D8601; end if; when s36AC7A0A1A83247FFEBA473A089671A1570A444F => if s38B47F4C3DE0DCB215428A00C075B72E81724995
 >= sE5CEEC534B45504250BB0AB9C68F528B4427B4EA then s1A1FBAC4E57E71A08D58F34D3F236E10FDBB13F1 <= '1'; if s42C156E01C093831B32D6A7CBFD3020F1F90D4CF = '1' then s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s3F5CD917DD715D35070C12A524859CBA336A5E8F; else s2A4FD558F206D02C009EE8C6C3270121218EBF72
 <= s4D060726C033C2FAEAF8BEA001EE62AE7781F8FF; end if; elsif s2352BDBE6CE03BBCE38F2DE675BB47F601C0CEE4 = '1' then s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s4E6FE1CA131098FC04443D071866EADE68B517F4; else s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s36AC7A0A1A83247FFEBA473A089671A1570A444F
; end if; when s4D060726C033C2FAEAF8BEA001EE62AE7781F8FF => if s38B47F4C3DE0DCB215428A00C075B72E81724995 >= sF1ACDF194238D93C80C3F56B982846A83ABF8042 then s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s4BD5B45FED6CFDC9C7C9EB134B11243E9E183FB8; elsif s2352BDBE6CE03BBCE38F2DE675BB47F601C0CEE4
 = '1' then s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s4E6FE1CA131098FC04443D071866EADE68B517F4; else s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s4D060726C033C2FAEAF8BEA001EE62AE7781F8FF; end if; when s4BD5B45FED6CFDC9C7C9EB134B11243E9E183FB8 => if s38B47F4C3DE0DCB215428A00C075B72E81724995
 >= s554B052BE2734AB000DFA8E34A6DCD1C5B7F62F3 then s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s3F5CD917DD715D35070C12A524859CBA336A5E8F; elsif s2352BDBE6CE03BBCE38F2DE675BB47F601C0CEE4 = '1' then s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s4E6FE1CA131098FC04443D071866EADE68B517F4
; else s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s4BD5B45FED6CFDC9C7C9EB134B11243E9E183FB8; end if; when s3F5CD917DD715D35070C12A524859CBA336A5E8F => if s38B47F4C3DE0DCB215428A00C075B72E81724995 >= sF18D65E9875B3783D0FD9B8A653B5F0B9BE8AE44 then s2A4FD558F206D02C009EE8C6C3270121218EBF72
 <= s39F04C15DE0E5F43C559F3657FACB1AA3D4A2CF7; elsif s2352BDBE6CE03BBCE38F2DE675BB47F601C0CEE4 = '1' then s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s4E6FE1CA131098FC04443D071866EADE68B517F4; else s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s3F5CD917DD715D35070C12A524859CBA336A5E8F
; end if; when s39F04C15DE0E5F43C559F3657FACB1AA3D4A2CF7 => if s803DC9CAA8B495BF1BF7AC678ABDB7265B406E97 = '1' and s45D2033B63004B619AF223745CE9944CA468D689 = '1' then s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= sC4E33B939FA9CAB7BA08E4FBF3DEF9689B5FB0C0;
 elsif s2352BDBE6CE03BBCE38F2DE675BB47F601C0CEE4 = '1' then s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s4E6FE1CA131098FC04443D071866EADE68B517F4; else s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s39F04C15DE0E5F43C559F3657FACB1AA3D4A2CF7; end if; when sC4E33B939FA9CAB7BA08E4FBF3DEF9689B5FB0C0
 => if s7BA0158498624EFFF7A85F2DE562B881D380F526 >= sA0F87C252F9449120B37FA8565AD3B246A3EBC17 then s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= sAC14180D3920A14E53EB388154EEB3BD8EE00F38; elsif s2352BDBE6CE03BBCE38F2DE675BB47F601C0CEE4 = '1' then s2A4FD558F206D02C009EE8C6C3270121218EBF72
 <= s4E6FE1CA131098FC04443D071866EADE68B517F4; else s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= sC4E33B939FA9CAB7BA08E4FBF3DEF9689B5FB0C0; end if; when sAC14180D3920A14E53EB388154EEB3BD8EE00F38 => if s7BA0158498624EFFF7A85F2DE562B881D380F526 >= s7D425144B574080EAE524904A8A3A1B003EE34A7
 then s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= sA265FC1FF568154C90487807499F4E4714E828D2; elsif s2352BDBE6CE03BBCE38F2DE675BB47F601C0CEE4 = '1' then s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s4E6FE1CA131098FC04443D071866EADE68B517F4; else s2A4FD558F206D02C009EE8C6C3270121218EBF72
 <= sAC14180D3920A14E53EB388154EEB3BD8EE00F38; end if; when sA265FC1FF568154C90487807499F4E4714E828D2 => if s7BA0158498624EFFF7A85F2DE562B881D380F526 >= s287FEDCA98AA2143D3F527A97C155CE0F210A782 then s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= sA8AD75438F0C3D62010B98FEDD21D5B11EF0BBC1
; elsif s2352BDBE6CE03BBCE38F2DE675BB47F601C0CEE4 = '1' then s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s4E6FE1CA131098FC04443D071866EADE68B517F4; else s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= sA265FC1FF568154C90487807499F4E4714E828D2; end if; when 
sA8AD75438F0C3D62010B98FEDD21D5B11EF0BBC1 => if s57AE96E3A4322EF36A1E1352A866E15B3C188F64='1' and s395EF2527A3109AD4086230A8FD7F23B1F2F0F41= '1' then s8DC239BAE0C4B59356AE3036500FFCCDBBFA8E72 <= '1'; s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s529B4ABD50A0DC309F792EE5D475A66D0D9959A2
; elsif s2352BDBE6CE03BBCE38F2DE675BB47F601C0CEE4 = '1' then s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s4E6FE1CA131098FC04443D071866EADE68B517F4; else s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= sA8AD75438F0C3D62010B98FEDD21D5B11EF0BBC1; end if; when 
s529B4ABD50A0DC309F792EE5D475A66D0D9959A2 => if s395EF2527A3109AD4086230A8FD7F23B1F2F0F41='0' then s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C; elsif s2352BDBE6CE03BBCE38F2DE675BB47F601C0CEE4 = '1' then s2A4FD558F206D02C009EE8C6C3270121218EBF72
 <= s4E6FE1CA131098FC04443D071866EADE68B517F4; else s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s529B4ABD50A0DC309F792EE5D475A66D0D9959A2; end if; when s4E6FE1CA131098FC04443D071866EADE68B517F4 =>  s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C
; when others => s2A4FD558F206D02C009EE8C6C3270121218EBF72 <= s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C; end case; end process s16A54A799612DE170F8EC9B0B99BAC7A233D1DF9;  s00506246AD19C23077849FB3ED52A1D57EAB8122 : process(clk_i) begin if rising_edge(clk_i
) then if reset_i = '1' then sEA8188CAD31707F17B299650F81C67D601FE09D7 <= (others => '0'); s2DE53BABF9E8291149A3F55C3450649370E3009F <= (others => '0'); sDF9F3E40D3B907510D4DF16BCDAFC2586EB30618 <= (others => '0'); s0465AAD501BCFB42A3CE710255F7BF6B54E619DD
 <= (others => '0'); s9216F1816ACE78FB0851459E9601420ABC3AA570 <= (others => '0'); s2C546333D09386C1C9D785047A9CEA69F8B26C94 <= (others => '0'); else  if s22E923CF436A1BF1EAA149BF66A7AD165ABABD9A=sBB12D33790A5D3018B4D986F4ADB83977C5D8601 then s0465AAD501BCFB42A3CE710255F7BF6B54E619DD
 <= (others => '0'); end if; if s22E923CF436A1BF1EAA149BF66A7AD165ABABD9A=s36AC7A0A1A83247FFEBA473A089671A1570A444F and s0FFAB4F8912FCE63B3997867066DFB9C1F628974='1' then sEA8188CAD31707F17B299650F81C67D601FE09D7 <= sEA8188CAD31707F17B299650F81C67D601FE09D7
(4 downto 0) & s395EF2527A3109AD4086230A8FD7F23B1F2F0F41; end if; if s22E923CF436A1BF1EAA149BF66A7AD165ABABD9A=s4D060726C033C2FAEAF8BEA001EE62AE7781F8FF and s0FFAB4F8912FCE63B3997867066DFB9C1F628974='1' then s2DE53BABF9E8291149A3F55C3450649370E3009F <= s2DE53BABF9E8291149A3F55C3450649370E3009F
(6 downto 0) & s395EF2527A3109AD4086230A8FD7F23B1F2F0F41; end if; if s22E923CF436A1BF1EAA149BF66A7AD165ABABD9A=s4BD5B45FED6CFDC9C7C9EB134B11243E9E183FB8 and s0FFAB4F8912FCE63B3997867066DFB9C1F628974='1' then sDF9F3E40D3B907510D4DF16BCDAFC2586EB30618 <= sDF9F3E40D3B907510D4DF16BCDAFC2586EB30618
(14 downto 0) & s395EF2527A3109AD4086230A8FD7F23B1F2F0F41; end if; if s22E923CF436A1BF1EAA149BF66A7AD165ABABD9A=sC4E33B939FA9CAB7BA08E4FBF3DEF9689B5FB0C0 and s45D2033B63004B619AF223745CE9944CA468D689='1' then s9216F1816ACE78FB0851459E9601420ABC3AA570(to_integer
(s7BA0158498624EFFF7A85F2DE562B881D380F526)) <= s395EF2527A3109AD4086230A8FD7F23B1F2F0F41; end if; if s22E923CF436A1BF1EAA149BF66A7AD165ABABD9A=sAC14180D3920A14E53EB388154EEB3BD8EE00F38 and s45D2033B63004B619AF223745CE9944CA468D689='1' then s0465AAD501BCFB42A3CE710255F7BF6B54E619DD
(to_integer(s7BA0158498624EFFF7A85F2DE562B881D380F526)) <= s395EF2527A3109AD4086230A8FD7F23B1F2F0F41; end if; if s22E923CF436A1BF1EAA149BF66A7AD165ABABD9A=sA265FC1FF568154C90487807499F4E4714E828D2 and s45D2033B63004B619AF223745CE9944CA468D689='1' then s2C546333D09386C1C9D785047A9CEA69F8B26C94
 <= s395EF2527A3109AD4086230A8FD7F23B1F2F0F41 & s2C546333D09386C1C9D785047A9CEA69F8B26C94(s2C546333D09386C1C9D785047A9CEA69F8B26C94'left downto 1); end if; end if; end if; end process s00506246AD19C23077849FB3ED52A1D57EAB8122; s08140CA014D79009968544D9ECD7EAA0E163EED4
 <= '1' when sEA8188CAD31707F17B299650F81C67D601FE09D7 = sD086456116C26514BAA46126BDD5342689EA4666 or sEA8188CAD31707F17B299650F81C67D601FE09D7 = s85EB2661C4F665AC828497B5A151BB556355E05B or  sEA8188CAD31707F17B299650F81C67D601FE09D7 = sAD320E17FE59D7A60E88C7BE1ADB0F57AA30EDD0
 or  sEA8188CAD31707F17B299650F81C67D601FE09D7 = sA4D53F04E8BA4766E83AD0DEFDD9278B52C3044C or  sEA8188CAD31707F17B299650F81C67D601FE09D7 = sEDFBFD9F8F54F1BD9B20E33D40221B2D6C287A4D or  sEA8188CAD31707F17B299650F81C67D601FE09D7 = s9B0C1672B259D9C1E1031A2B01F0DF6FE98F2A2E
 or  sEA8188CAD31707F17B299650F81C67D601FE09D7 = sE78665F3E53F7F72C28BF19FCA20946AD4B10D08 else  '0'; s7D425144B574080EAE524904A8A3A1B003EE34A7 <= to_unsigned(sF073296EFBB46BD30ADC8EA25E1CC93687EBDAFB,32) when sEA8188CAD31707F17B299650F81C67D601FE09D7 = sD086456116C26514BAA46126BDD5342689EA4666
 or sEA8188CAD31707F17B299650F81C67D601FE09D7 = s85EB2661C4F665AC828497B5A151BB556355E05B or sEA8188CAD31707F17B299650F81C67D601FE09D7 = sAD320E17FE59D7A60E88C7BE1ADB0F57AA30EDD0 or sEA8188CAD31707F17B299650F81C67D601FE09D7 = sA4D53F04E8BA4766E83AD0DEFDD9278B52C3044C
 or sEA8188CAD31707F17B299650F81C67D601FE09D7 = sEDFBFD9F8F54F1BD9B20E33D40221B2D6C287A4D or  sEA8188CAD31707F17B299650F81C67D601FE09D7 = s9B0C1672B259D9C1E1031A2B01F0DF6FE98F2A2E or sEA8188CAD31707F17B299650F81C67D601FE09D7 = sE78665F3E53F7F72C28BF19FCA20946AD4B10D08
 else to_unsigned(41,32) when sEA8188CAD31707F17B299650F81C67D601FE09D7 = sA2C6EE455D0B31BBD6DC87409C4BCCEE5CFD35BD else to_unsigned(24,32);  sA0F87C252F9449120B37FA8565AD3B246A3EBC17 <= x"00000000" when sEA8188CAD31707F17B299650F81C67D601FE09D7 = sC950D600C869099649CD1A85609BA2714F805E57
 or sEA8188CAD31707F17B299650F81C67D601FE09D7 = s37EC8A8DDC24DE5CCA325C6D520F09FE8B8BE3B0 or  sEA8188CAD31707F17B299650F81C67D601FE09D7 = sCE667A08F3FDC358AF7C3578CD6983F0DD93374C or  sEA8188CAD31707F17B299650F81C67D601FE09D7 = sEFA6395FD066E102662C9126CF88821C4940A5E2
 or  sEA8188CAD31707F17B299650F81C67D601FE09D7 = sA2C6EE455D0B31BBD6DC87409C4BCCEE5CFD35BD or  sEA8188CAD31707F17B299650F81C67D601FE09D7 = sBB116EDD54150FE461AF440792906CBAF166BCC9 else  x"00000001" when sEA8188CAD31707F17B299650F81C67D601FE09D7 = sD086456116C26514BAA46126BDD5342689EA4666
 else x"00000002" when sEA8188CAD31707F17B299650F81C67D601FE09D7 = s85EB2661C4F665AC828497B5A151BB556355E05B or sEA8188CAD31707F17B299650F81C67D601FE09D7 = sAD320E17FE59D7A60E88C7BE1ADB0F57AA30EDD0 or sEA8188CAD31707F17B299650F81C67D601FE09D7 = sA4D53F04E8BA4766E83AD0DEFDD9278B52C3044C
 or sEA8188CAD31707F17B299650F81C67D601FE09D7 = sEDFBFD9F8F54F1BD9B20E33D40221B2D6C287A4D or sEA8188CAD31707F17B299650F81C67D601FE09D7 = s9B0C1672B259D9C1E1031A2B01F0DF6FE98F2A2E or sEA8188CAD31707F17B299650F81C67D601FE09D7 = sE78665F3E53F7F72C28BF19FCA20946AD4B10D08
 else x"00000000";   s42C156E01C093831B32D6A7CBFD3020F1F90D4CF <= '0' when sEA8188CAD31707F17B299650F81C67D601FE09D7 = sC950D600C869099649CD1A85609BA2714F805E57 or sEA8188CAD31707F17B299650F81C67D601FE09D7 = s37EC8A8DDC24DE5CCA325C6D520F09FE8B8BE3B0 or sEA8188CAD31707F17B299650F81C67D601FE09D7
 = sCE667A08F3FDC358AF7C3578CD6983F0DD93374C or sEA8188CAD31707F17B299650F81C67D601FE09D7 = sEFA6395FD066E102662C9126CF88821C4940A5E2 or sEA8188CAD31707F17B299650F81C67D601FE09D7 = s01C3860AF9A5F5F7A28F043ECA30EAB1DE4D786E or sEA8188CAD31707F17B299650F81C67D601FE09D7
 = sA2C6EE455D0B31BBD6DC87409C4BCCEE5CFD35BD else '1';  s22BF2481500BFBC968E4E77572AF70B5D2314799 : process(clk_i) begin if rising_edge(clk_i) then if reset_i='1' then s38B47F4C3DE0DCB215428A00C075B72E81724995 <= (others => '0'); else if s22E923CF436A1BF1EAA149BF66A7AD165ABABD9A
 /= s2A4FD558F206D02C009EE8C6C3270121218EBF72 then s38B47F4C3DE0DCB215428A00C075B72E81724995 <= (others => '0'); elsif s0FFAB4F8912FCE63B3997867066DFB9C1F628974='1' then s38B47F4C3DE0DCB215428A00C075B72E81724995 <= s38B47F4C3DE0DCB215428A00C075B72E81724995
 + 1; end if; end if; end if; end process s22BF2481500BFBC968E4E77572AF70B5D2314799; s11F5C144354B941A399EDCA7F8F883E698605F11 : process(clk_i) begin if rising_edge(clk_i) then if reset_i='1' then sDEB77204C753BE668599CE98F2768D24342B4D6B <= '0'; else sDEB77204C753BE668599CE98F2768D24342B4D6B
 <= s44987DF76FE68D9CEF103968757796A160C63E1C; end if; end if; end process s11F5C144354B941A399EDCA7F8F883E698605F11; s44987DF76FE68D9CEF103968757796A160C63E1C <= '1' when s2A4FD558F206D02C009EE8C6C3270121218EBF72 = s39F04C15DE0E5F43C559F3657FACB1AA3D4A2CF7
 and s22E923CF436A1BF1EAA149BF66A7AD165ABABD9A /= s39F04C15DE0E5F43C559F3657FACB1AA3D4A2CF7 else  '0' when s1E9AD3357247BE14ACDD8BA1FE752CC280C75D49 = '1' else  sDEB77204C753BE668599CE98F2768D24342B4D6B; s63964CD9864321E03FA6345CE209189BDF142292 : process
(clk_i) begin if rising_edge(clk_i) then if reset_i='1' then s803DC9CAA8B495BF1BF7AC678ABDB7265B406E97 <= '0'; else s803DC9CAA8B495BF1BF7AC678ABDB7265B406E97 <= s8E9F68EAF8B9CC6752ACCB89FC9C7B7337F6BBA7; end if; end if; end process s63964CD9864321E03FA6345CE209189BDF142292
; s8E9F68EAF8B9CC6752ACCB89FC9C7B7337F6BBA7 <= '1' when s1E9AD3357247BE14ACDD8BA1FE752CC280C75D49 = '1' else  '0' when s2A4FD558F206D02C009EE8C6C3270121218EBF72 = s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C else  s803DC9CAA8B495BF1BF7AC678ABDB7265B406E97;  
s18EE0CA54CE5DCA3FF51E54A534422E5289F2878 : process(clk_i) begin if rising_edge(clk_i) then if reset_i='1' then s9E27824C43FC3BC94286CC02E57D7EA018AB2D12 <= (others => '0'); elsif sDEB77204C753BE668599CE98F2768D24342B4D6B = '1' then if s0FFAB4F8912FCE63B3997867066DFB9C1F628974
='1' then s9E27824C43FC3BC94286CC02E57D7EA018AB2D12 <= (others => '0'); elsif s9E27824C43FC3BC94286CC02E57D7EA018AB2D12 < 127 then s9E27824C43FC3BC94286CC02E57D7EA018AB2D12 <= s9E27824C43FC3BC94286CC02E57D7EA018AB2D12 + 1; end if; end if; end if; end process
 s18EE0CA54CE5DCA3FF51E54A534422E5289F2878; s1E9AD3357247BE14ACDD8BA1FE752CC280C75D49 <= '1' when sDEB77204C753BE668599CE98F2768D24342B4D6B='1' and (s395EF2527A3109AD4086230A8FD7F23B1F2F0F41 = '0' and sC3ADFA536EF4E4699F020FEC7F3F5E5F95645E71 = '1') else '0';
  s88F91B1F3C95788B28B86AFE7AF74EAE6DE03121 : process(clk_i) begin if rising_edge(clk_i) then if reset_i='1' then sA2DAE05A577AC12D23A3CED89B449A366DCFF9D3 <= (others => '0'); s5960FAE099FE1D30E1893ED128A9BC168134F816 <= '0'; elsif s5960FAE099FE1D30E1893ED128A9BC168134F816
 = '0' then if s1E9AD3357247BE14ACDD8BA1FE752CC280C75D49 = '1' then sA2DAE05A577AC12D23A3CED89B449A366DCFF9D3 <= s9E27824C43FC3BC94286CC02E57D7EA018AB2D12; s5960FAE099FE1D30E1893ED128A9BC168134F816 <= '1'; end if; end if; end if; end process s88F91B1F3C95788B28B86AFE7AF74EAE6DE03121
; s5F9BC299EFE239681824EDA47F57D2770C69A4E4 : process(clk_i) begin if rising_edge(clk_i) then if reset_i='1' then s7BA0158498624EFFF7A85F2DE562B881D380F526 <= (others => '0'); elsif s22E923CF436A1BF1EAA149BF66A7AD165ABABD9A /= s2A4FD558F206D02C009EE8C6C3270121218EBF72
 then s7BA0158498624EFFF7A85F2DE562B881D380F526 <= (others => '0'); elsif s45D2033B63004B619AF223745CE9944CA468D689='1' then s7BA0158498624EFFF7A85F2DE562B881D380F526 <= s7BA0158498624EFFF7A85F2DE562B881D380F526 + 1; end if; end if; end process s5F9BC299EFE239681824EDA47F57D2770C69A4E4
;  s5D5A3E73528088194AE8DEF5C45CAE334B300752 : process(clk_i) begin if rising_edge(clk_i) then if reset_i='1' then s299A4649AF76D252E8BCE9B9976634617E034DC3 <= (others => '0'); else if s22E923CF436A1BF1EAA149BF66A7AD165ABABD9A /= s2A4FD558F206D02C009EE8C6C3270121218EBF72
 then s299A4649AF76D252E8BCE9B9976634617E034DC3 <= (others => '0'); else s299A4649AF76D252E8BCE9B9976634617E034DC3 <= s299A4649AF76D252E8BCE9B9976634617E034DC3 + 1; end if; end if; end if; end process s5D5A3E73528088194AE8DEF5C45CAE334B300752;   s2BC74474AF6817AD93D4AB843A4D19F0B6E381AD
 : process(clk_i) begin if rising_edge(clk_i) then if reset_i='1' then s2F285CF0B57A3B502B36C687EFD83233AC8934DC <= (others => '0'); else if s57AE96E3A4322EF36A1E1352A866E15B3C188F64='0' then s2F285CF0B57A3B502B36C687EFD83233AC8934DC <= (others => '0'); elsif
 s2F285CF0B57A3B502B36C687EFD83233AC8934DC < unsigned(tReset_i) then s2F285CF0B57A3B502B36C687EFD83233AC8934DC <= s2F285CF0B57A3B502B36C687EFD83233AC8934DC + 1; end if; end if; end if; end process s2BC74474AF6817AD93D4AB843A4D19F0B6E381AD; s2352BDBE6CE03BBCE38F2DE675BB47F601C0CEE4
 <= '1' when s2F285CF0B57A3B502B36C687EFD83233AC8934DC >= unsigned(tReset_i) else '0';  sF073296EFBB46BD30ADC8EA25E1CC93687EBDAFB <= to_integer(unsigned(numPulPosVal_i));    s1ECA68304446F3295D7FC3C5B314ADBA0067C044 <= to_integer(unsigned(distRev_i)); sB3A8B19CA98570BA8D1B96F098A8058070AA0E06
 <= to_integer(unsigned(numPulPosVal_i)); s495F0760A6D370CF2E5DACC3A884F77824629006 : process(sB3A8B19CA98570BA8D1B96F098A8058070AA0E06, s0465AAD501BCFB42A3CE710255F7BF6B54E619DD, sEA8188CAD31707F17B299650F81C67D601FE09D7, s1ECA68304446F3295D7FC3C5B314ADBA0067C044
) begin  s38FBA08FA1E8936955F6D21A792256E3658F8387 <= (others => '0'); s6D8E140706515F7AFC288159A5BC35A838C23C32 <= (others => '0'); case sEA8188CAD31707F17B299650F81C67D601FE09D7 is when sD086456116C26514BAA46126BDD5342689EA4666 | s85EB2661C4F665AC828497B5A151BB556355E05B
 | sAD320E17FE59D7A60E88C7BE1ADB0F57AA30EDD0 | sA4D53F04E8BA4766E83AD0DEFDD9278B52C3044C | sEDFBFD9F8F54F1BD9B20E33D40221B2D6C287A4D | s9B0C1672B259D9C1E1031A2B01F0DF6FE98F2A2E | sE78665F3E53F7F72C28BF19FCA20946AD4B10D08 => for s020F5125771EEEB6F963720A8BB968FCA977AA41
 in 0 to 31 loop if (s020F5125771EEEB6F963720A8BB968FCA977AA41 < s1ECA68304446F3295D7FC3C5B314ADBA0067C044) then s6D8E140706515F7AFC288159A5BC35A838C23C32(s020F5125771EEEB6F963720A8BB968FCA977AA41) <= s0465AAD501BCFB42A3CE710255F7BF6B54E619DD(s020F5125771EEEB6F963720A8BB968FCA977AA41
 + (sB3A8B19CA98570BA8D1B96F098A8058070AA0E06-s1ECA68304446F3295D7FC3C5B314ADBA0067C044)); end if; if (s020F5125771EEEB6F963720A8BB968FCA977AA41 < sB3A8B19CA98570BA8D1B96F098A8058070AA0E06-s1ECA68304446F3295D7FC3C5B314ADBA0067C044) then s38FBA08FA1E8936955F6D21A792256E3658F8387
(s020F5125771EEEB6F963720A8BB968FCA977AA41) <= s0465AAD501BCFB42A3CE710255F7BF6B54E619DD(s020F5125771EEEB6F963720A8BB968FCA977AA41); end if; end loop; when sCE667A08F3FDC358AF7C3578CD6983F0DD93374C | sC950D600C869099649CD1A85609BA2714F805E57 | s37EC8A8DDC24DE5CCA325C6D520F09FE8B8BE3B0
 | sEFA6395FD066E102662C9126CF88821C4940A5E2 | s01C3860AF9A5F5F7A28F043ECA30EAB1DE4D786E | sBB116EDD54150FE461AF440792906CBAF166BCC9 => s38FBA08FA1E8936955F6D21A792256E3658F8387(15 downto 0) <= s0465AAD501BCFB42A3CE710255F7BF6B54E619DD(15 downto 0); s6D8E140706515F7AFC288159A5BC35A838C23C32
 <= (others => '0'); when sA2C6EE455D0B31BBD6DC87409C4BCCEE5CFD35BD =>  s38FBA08FA1E8936955F6D21A792256E3658F8387(31 downto 0) <= s0465AAD501BCFB42A3CE710255F7BF6B54E619DD(31 downto 0); s6D8E140706515F7AFC288159A5BC35A838C23C32(7 downto 0) <= s0465AAD501BCFB42A3CE710255F7BF6B54E619DD
(39 downto 32); when others => s38FBA08FA1E8936955F6D21A792256E3658F8387 <= (others => '0'); s6D8E140706515F7AFC288159A5BC35A838C23C32 <= (others => '0'); end case; end process s495F0760A6D370CF2E5DACC3A884F77824629006;  s4F8EEACE44418C026D8F7B6609F95D9F2983F61C
 <= s9216F1816ACE78FB0851459E9601420ABC3AA570(0); sEB2C0A31F86ED13FF0CDECB77CA291A86128B247 <= s9216F1816ACE78FB0851459E9601420ABC3AA570(1);    s98683DAEF246D4975C386EA22C561360083D1221 : process(clk_i) begin if rising_edge(clk_i) then if reset_i = '1' then
 dataValid_o <= '0'; rxPosVal_o <= (others => '0'); numRev_o <= (others => '0'); error_o <= (others => '0'); else  dataValid_o <= '0';  if s8DC239BAE0C4B59356AE3036500FFCCDBBFA8E72='1' and s08140CA014D79009968544D9ECD7EAA0E163EED4='1' then rxPosVal_o <= s38FBA08FA1E8936955F6D21A792256E3658F8387
; numRev_o <= s6D8E140706515F7AFC288159A5BC35A838C23C32;  end if;  if s22E923CF436A1BF1EAA149BF66A7AD165ABABD9A = s529B4ABD50A0DC309F792EE5D475A66D0D9959A2 and s2A4FD558F206D02C009EE8C6C3270121218EBF72 = s2AAC85453BFE1F0ECA7CE3219C0D858541D7495C and s08140CA014D79009968544D9ECD7EAA0E163EED4
='1' then dataValid_o <= '1'; end if; end if; end if; end process s98683DAEF246D4975C386EA22C561360083D1221; end struct;