library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;
  
  use work.BISS_pkg.all;

entity BISS is
  port
  (
    clk_i             : in std_logic;
    reset_i           : in std_logic;
    
    version           : out std_logic_vector(31 downto 0);     
    
    clockDiv_i        : in std_logic_vector(31 downto 0);
    startCmd_i        : in std_logic;                     
    numBits_i         : in std_logic_vector(7 downto 0);  
    timeOutClkCount_i : in std_logic_vector (15 downto 0);   
    
    dataRxWord01_o    : out std_logic_vector(31 downto 0);
    dataRxWord02_o    : out std_logic_vector(31 downto 0);
    dataValid_o       : out std_logic;      
    error_o           : out std_logic;
    
    MA_o              : out std_logic;
    SLI_i             : in  std_logic;
    SLO_o             : out std_logic 
  );
end BISS;

architecture struct OF BISS IS  signal s6B30F3AB3E2DD07A9ECE5389D13080965A495139 : std_logic_vector(63 downto 0); signal sD81661E305E822B9113FF02F9996CA02905AC938 : std_logic; signal s04275C0AE3DFB7E3AC35D244C846CE3E529EAF44 : std_logic; signal s260631C53159B3E5FCFC9E4888313F57276113A3
 : std_logic; signal s3A269885069B7EEA657EF3DED6121E17648A8490 : std_logic; signal s46ABF5D9FEA69A802E945C6413E9BEF020D86842 : std_logic; begin version <= "10" & s731A256AA7EC109FE962BF102445534C5772925D & s7EC4167F3F7F1E99D074313BF18FF4BA05E7ED10 & s5907A17D8E29C7EB61D4F347241BFE4DAC407AEA
;    s6BD109C578CF89126A14BF943E8522A9004A7540: entity work.BISS_clockGen port map ( s82C78E3CD667612DE97ED7C5FA8365F21045093F => clk_i, s0A61EC3B284D41A7527B973B71395AF396BD0749 => reset_i, s1C654E69626584446DE718F7EE7988BA2A365CCF => clockDiv_i, s36AD3DDD0D7E89B06FC50291B7727A74872462C3
 => sD81661E305E822B9113FF02F9996CA02905AC938, s1FDEC574EB5E12EA0B4DDD4FCA57414E037CB358 => s04275C0AE3DFB7E3AC35D244C846CE3E529EAF44,  s35446BFB0A5C8D55EEA546BF7816F1ECD3A67612 => s260631C53159B3E5FCFC9E4888313F57276113A3, s011A91380BC90B6ACF14422413DCD2C29E155965
 => s3A269885069B7EEA657EF3DED6121E17648A8490, sDC4EF638ACF00C773A1E6DC2D7F59B1ED9BE8A9F => s46ABF5D9FEA69A802E945C6413E9BEF020D86842 ); s2373A2787FACCE2B357A5B86FA3FEAEA1748C512: entity work.BISS_control port map ( s82C78E3CD667612DE97ED7C5FA8365F21045093F
 => clk_i, s0A61EC3B284D41A7527B973B71395AF396BD0749 => reset_i, sEC9D498A27032D5D5CC9FBE9786A936DA84A5766 => s3A269885069B7EEA657EF3DED6121E17648A8490, sADBC8E7E04FA85F5322F3AAA6BF0398152DF9E93 => s46ABF5D9FEA69A802E945C6413E9BEF020D86842, s67AA1F47031AD081937F209C8CEB3917E3285B98
 => startCmd_i, sBF63B84FE256F013F6F36AB8B222082B8647B811 => numBits_i, s865C7DE113F62D5D7CAC52C2E96B9519EB8FF306 => timeOutClkCount_i, sE9D5A330018FD42F21BED92AE3F25BEBD3119C81 => sD81661E305E822B9113FF02F9996CA02905AC938, s8D52A510B7F21BBB60B0674B11C3DA67D5DE5713
 => s04275C0AE3DFB7E3AC35D244C846CE3E529EAF44, s6C6651D383B41FAFDF50F2BAA251FDC2A08AB191 => dataValid_o, s4F8467F3FA446F57411E855E04FB8C5F7C144A28 => s6B30F3AB3E2DD07A9ECE5389D13080965A495139, sE4ED7921C578950CCEB828999E51D6DAE12F5A90 => error_o,  s4088069AAB16D293A7469FD360A0287D49DE79AE
 => s260631C53159B3E5FCFC9E4888313F57276113A3, s76D10F4B556F2B64C06E85300CE7EC78B730048A => SLI_i );  dataRxWord01_o <= s6B30F3AB3E2DD07A9ECE5389D13080965A495139( 31 downto 0); dataRxWord02_o <= s6B30F3AB3E2DD07A9ECE5389D13080965A495139( 63 downto 32); MA_o
 <= s260631C53159B3E5FCFC9E4888313F57276113A3; SLO_o <= '0'; end struct;