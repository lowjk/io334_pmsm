library ieee; use ieee.std_logic_1164.all; use ieee.numeric_std.all; entity BISS_clockGen is port ( s82C78E3CD667612DE97ED7C5FA8365F21045093F : in std_logic; s0A61EC3B284D41A7527B973B71395AF396BD0749 : in std_logic; s1C654E69626584446DE718F7EE7988BA2A365CCF
 : in std_logic_vector(31 downto 0); s36AD3DDD0D7E89B06FC50291B7727A74872462C3 : in std_logic; s1FDEC574EB5E12EA0B4DDD4FCA57414E037CB358 : in std_logic;  s35446BFB0A5C8D55EEA546BF7816F1ECD3A67612 : out std_logic; s011A91380BC90B6ACF14422413DCD2C29E155965 : 
out std_logic; sDC4EF638ACF00C773A1E6DC2D7F59B1ED9BE8A9F : out std_logic ); end BISS_clockGen; architecture rtl of BISS_clockGen is type s7F0B6A4643B458243E2E60698CD8F724E1B5692D is (s03D0DCDB162423DE6D6DEA3D2A6DCAEEBE3FAE63, s3B85CA1896C05344D1B0F452D7CF00D8590562E3
, sC02F7EF233036620CCCD2F33AA9C747216F23696); signal s1C8654799AD97A5646787FCC52F12F0D731697D9, s5B32DB06E10FB9324A8A8C8CADE6A1B29B288A8E : s7F0B6A4643B458243E2E60698CD8F724E1B5692D; signal s260631C53159B3E5FCFC9E4888313F57276113A3 : std_logic; signal s2CC9648F3BE766AD963F4674275246BB5BDC578E
 : std_logic; signal s38B47F4C3DE0DCB215428A00C075B72E81724995 : unsigned(31 downto 0); signal s3D815B08D1A39BF5E3E1B838DF0F21DA44D5A015 : std_logic; signal s31AFBA8FA30A69D2BF8C4A74E99AF3A6667AB1BB : std_logic; begin s1B8DE4320EEAE9B0C4ABE0C0EAA1B6335C6FE6C8
: process(s1C8654799AD97A5646787FCC52F12F0D731697D9, s36AD3DDD0D7E89B06FC50291B7727A74872462C3, s1FDEC574EB5E12EA0B4DDD4FCA57414E037CB358, s1C654E69626584446DE718F7EE7988BA2A365CCF, s38B47F4C3DE0DCB215428A00C075B72E81724995) begin  s260631C53159B3E5FCFC9E4888313F57276113A3
 <= '1'; case s1C8654799AD97A5646787FCC52F12F0D731697D9 is when s03D0DCDB162423DE6D6DEA3D2A6DCAEEBE3FAE63 => s260631C53159B3E5FCFC9E4888313F57276113A3 <= '1'; if s36AD3DDD0D7E89B06FC50291B7727A74872462C3='1' then s5B32DB06E10FB9324A8A8C8CADE6A1B29B288A8E <= 
s3B85CA1896C05344D1B0F452D7CF00D8590562E3; else s5B32DB06E10FB9324A8A8C8CADE6A1B29B288A8E <= s03D0DCDB162423DE6D6DEA3D2A6DCAEEBE3FAE63; end if; when s3B85CA1896C05344D1B0F452D7CF00D8590562E3 => s260631C53159B3E5FCFC9E4888313F57276113A3 <= '0'; if s1FDEC574EB5E12EA0B4DDD4FCA57414E037CB358
='1' then s5B32DB06E10FB9324A8A8C8CADE6A1B29B288A8E <= s03D0DCDB162423DE6D6DEA3D2A6DCAEEBE3FAE63; elsif s38B47F4C3DE0DCB215428A00C075B72E81724995 >= unsigned(s1C654E69626584446DE718F7EE7988BA2A365CCF)-1 then s5B32DB06E10FB9324A8A8C8CADE6A1B29B288A8E <= sC02F7EF233036620CCCD2F33AA9C747216F23696
; else s5B32DB06E10FB9324A8A8C8CADE6A1B29B288A8E <= s3B85CA1896C05344D1B0F452D7CF00D8590562E3; end if; when sC02F7EF233036620CCCD2F33AA9C747216F23696 => s260631C53159B3E5FCFC9E4888313F57276113A3 <= '1'; if s1FDEC574EB5E12EA0B4DDD4FCA57414E037CB358='1' then
 s5B32DB06E10FB9324A8A8C8CADE6A1B29B288A8E <= s03D0DCDB162423DE6D6DEA3D2A6DCAEEBE3FAE63; elsif s38B47F4C3DE0DCB215428A00C075B72E81724995 >= unsigned(s1C654E69626584446DE718F7EE7988BA2A365CCF)-1 then s5B32DB06E10FB9324A8A8C8CADE6A1B29B288A8E <= s3B85CA1896C05344D1B0F452D7CF00D8590562E3
; else s5B32DB06E10FB9324A8A8C8CADE6A1B29B288A8E <= sC02F7EF233036620CCCD2F33AA9C747216F23696; end if; end case; end process s1B8DE4320EEAE9B0C4ABE0C0EAA1B6335C6FE6C8;  s01B836CC599AAC170C41C635FD46B72FA2B88119: process(s82C78E3CD667612DE97ED7C5FA8365F21045093F
, s0A61EC3B284D41A7527B973B71395AF396BD0749) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749 = '1' then s1C8654799AD97A5646787FCC52F12F0D731697D9 <= s03D0DCDB162423DE6D6DEA3D2A6DCAEEBE3FAE63; elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) 
then s1C8654799AD97A5646787FCC52F12F0D731697D9 <= s5B32DB06E10FB9324A8A8C8CADE6A1B29B288A8E; end if; end process s01B836CC599AAC170C41C635FD46B72FA2B88119;  s80E6945E63F32295F00E21A70F3B1647AFED9E48 : process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749
) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749='1' then s38B47F4C3DE0DCB215428A00C075B72E81724995 <= (others => '0'); elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then if s1C8654799AD97A5646787FCC52F12F0D731697D9 /= s5B32DB06E10FB9324A8A8C8CADE6A1B29B288A8E
 then s38B47F4C3DE0DCB215428A00C075B72E81724995 <= (others => '0'); else s38B47F4C3DE0DCB215428A00C075B72E81724995 <= s38B47F4C3DE0DCB215428A00C075B72E81724995 + 1; end if; end if; end process s80E6945E63F32295F00E21A70F3B1647AFED9E48;  s1DDD5F0829B5CE25CBF9A343410FB0DA516D24D6
: process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749='1' then s2CC9648F3BE766AD963F4674275246BB5BDC578E <= '0'; elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F
) then s2CC9648F3BE766AD963F4674275246BB5BDC578E <= s260631C53159B3E5FCFC9E4888313F57276113A3; end if; end process s1DDD5F0829B5CE25CBF9A343410FB0DA516D24D6; s3D815B08D1A39BF5E3E1B838DF0F21DA44D5A015 <= '1' when s2CC9648F3BE766AD963F4674275246BB5BDC578E='0' 
and s260631C53159B3E5FCFC9E4888313F57276113A3='1' else '0'; s31AFBA8FA30A69D2BF8C4A74E99AF3A6667AB1BB <= '1' when s2CC9648F3BE766AD963F4674275246BB5BDC578E='1' and s260631C53159B3E5FCFC9E4888313F57276113A3='0' else '0';  s35446BFB0A5C8D55EEA546BF7816F1ECD3A67612
 <= s260631C53159B3E5FCFC9E4888313F57276113A3; s011A91380BC90B6ACF14422413DCD2C29E155965 <= s3D815B08D1A39BF5E3E1B838DF0F21DA44D5A015; sDC4EF638ACF00C773A1E6DC2D7F59B1ED9BE8A9F <= s31AFBA8FA30A69D2BF8C4A74E99AF3A6667AB1BB; end rtl;