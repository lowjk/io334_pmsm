library IEEE; use IEEE.STD_LOGIC_1164.ALL; use IEEE.Numeric_Std.all; entity QAE_POSITIONNER is port( s2BE12327C739923A0BDA5AD372381D3F992B6A0F : in std_logic_vector(31 downto 0); s90724AE20811A4A1CF4892AD6C5DE35913A379E1 : in std_logic; s8EC1CD656701F1799C089F63518E2F895FE6470D
 : in std_logic; sDF13852084C1BE285B56723469BE3ADFFCF3653B : in std_logic_vector(31 downto 0); sE3594CA1813735566777C0F293E54987EE6AC901 : out std_logic ); end QAE_POSITIONNER; architecture rtl of QAE_POSITIONNER is begin sE3594CA1813735566777C0F293E54987EE6AC901
 <= '1' when s90724AE20811A4A1CF4892AD6C5DE35913A379E1 = '1' and s8EC1CD656701F1799C089F63518E2F895FE6470D = '1' else '1' when s90724AE20811A4A1CF4892AD6C5DE35913A379E1 = '1' and sDF13852084C1BE285B56723469BE3ADFFCF3653B /= s2BE12327C739923A0BDA5AD372381D3F992B6A0F
 and s8EC1CD656701F1799C089F63518E2F895FE6470D = '0' else '0'; end rtl; 