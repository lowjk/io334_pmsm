library ieee; use ieee.std_logic_1164.all; package BISS_ENCODER_pkg is  constant s731A256AA7EC109FE962BF102445534C5772925D : std_logic_vector(9 DOWNTO 0) := "00" & x"12";  constant s7EC4167F3F7F1E99D074313BF18FF4BA05E7ED10 : std_logic_vector(9 DOWNTO 0) := "00" & x"01";
 constant s5907A17D8E29C7EB61D4F347241BFE4DAC407AEA : std_logic_vector(9 DOWNTO 0) := "00" & x"06"; end BISS_ENCODER_pkg; 