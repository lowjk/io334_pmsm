library ieee; use ieee.std_logic_1164.all; package ENDAT_ENCODER_pkg is  constant s731A256AA7EC109FE962BF102445534C5772925D : std_logic_vector(9 DOWNTO 0) := "00" & x"1A";  constant s7EC4167F3F7F1E99D074313BF18FF4BA05E7ED10 : std_logic_vector(9 DOWNTO 0) := "00" & x"01";
 constant s5907A17D8E29C7EB61D4F347241BFE4DAC407AEA : std_logic_vector(9 DOWNTO 0) := "00" & x"02";    constant sDAD1E1924BFE7487D5AA58FB0E3AB6D80AFF7D81 : integer:= 6;  constant s8C1FCFB0787BDC32C8C8E0A79092BFBF8C9B3B95 : integer:= 7;  constant s2B661762AEA08905D55D9C993A5A3B37FF2EC6CD
 : integer:= 32;  constant sCD3268FB2E69A058B357988C1BAD31C26B18C0D3 : integer:= 56;   constant s1E05517C0679F267FA88812F99D44A02FF4ED0F5 : std_logic_vector(5 downto 0) := "000111";  constant sB64238E7DDBD6F205572B1E9360AE1265D8B4AEA : std_logic_vector(5 
downto 0) := "001110";  constant s3CE74FA91201742DE9903A95D23643FE5849757A : std_logic_vector(5 downto 0) := "010101";  constant s577F58458D046FA77A685C62ED8B8FEF8CDC09C9 : std_logic_vector(5 downto 0) := "011100";  constant s552E31DD6EF995EED1A8B6C12E49DC2C0A51F02F
 : std_logic_vector(5 downto 0) := "100011";  constant sFD1F530F2A18F9FF75CACE3E3D4051529EEF6982 : std_logic_vector(5 downto 0) := "101010";  constant s4BAA4FCE531A4298A40EF2ED066D556B6C1ECA42 : std_logic_vector(5 downto 0) := "110001";  constant s6DF2D092E032E7162C3A0DCC2D5A97E7D64555CC
 : std_logic_vector(5 downto 0) := "111000";  constant s7C44A19C549366606448A233C29ACDE5E6A81157 : std_logic_vector(5 downto 0) := "001001";  constant sC8DFB6E167EC00F6006ED436F19C33DEA279EBB8 : std_logic_vector(5 downto 0) := "010010";  constant s1BBF2B23FDB75A9E9E9C8410C6BD529018F0523E
 : std_logic_vector(5 downto 0) := "011011";  constant s57B57A47070F7BCB8EEBBEEA644F26DD6561AA10 : std_logic_vector(5 downto 0) := "100100";  constant sEF8743F14736EEC37C81CB3F1D2B016A785A0472 : std_logic_vector(5 downto 0) := "101101";  constant s467E7002675271D0D9C72D30C95CAD20E650A403
 : std_logic_vector(5 downto 0) := "110110";   constant sC467071B4163DF3B730A3D8FDBA24B62A24337A7 : std_logic_vector(7 downto 0) := x"40"; constant s497A41403D0E1204014E9B612AD737C8D35B3826 : std_logic_vector(7 downto 0) := x"41"; constant sFA0C0FC5DB4F0920FD931E78C8F3FFB13715D3FD
 : std_logic_vector(7 downto 0) := x"42"; constant s0E620B5ED6FCC4C01B20B593ADCB3709FA0BE26E : std_logic_vector(7 downto 0) := x"43"; constant s5AE40AED79A09E5B98B32D981F056406C9D6D977 : std_logic_vector(7 downto 0) := x"44"; constant sF76D4DB16EF1ADE5770C213F52561503D34DEF48
 : std_logic_vector(7 downto 0) := x"45"; constant sFE54C7D0CC6A2E8CFA4216501DCE1D8F436FEDC6 : std_logic_vector(7 downto 0) := x"46"; constant s7840E41D30357FC6180671D694922360D68CC896 : std_logic_vector(7 downto 0) := x"47"; constant sB8FBD8D6BBEDF46E31A0507EABC8F686CFB5CFA0
 : std_logic_vector(7 downto 0) := x"48"; constant s41500258240C5111284D79C684750BDFCF9BB4C9 : std_logic_vector(7 downto 0) := x"49"; constant s726B1776BF9E9357377F4BD979D5C542A12D7ECE : std_logic_vector(7 downto 0) := x"4A"; constant s83ADFBE2A97ACC106909DAC843AFC39378B31F29
 : std_logic_vector(7 downto 0) := x"4B"; constant sCF680DC8F214E3DEE1C42E950A30559BBAC4F3EB : std_logic_vector(7 downto 0) := x"4C"; constant s030F867793634A136982960F35AEAEFADF3FF2E0 : std_logic_vector(7 downto 0) := x"4D"; constant sDB159321904E6E9F130985F9B9AA585A8C6A0047
 : std_logic_vector(7 downto 0) := x"4E"; constant s57E60BF34E25CCC564142C57DBFF63876615DB5E : std_logic_vector(7 downto 0) := x"4F";  constant s190163C428AF25FC3187CA8FA8195F66129DEE18 : std_logic_vector(7 downto 0) := x"50"; constant sD753454CEAEA82A91076ECB6EF4A5F2112BC34A0
 : std_logic_vector(7 downto 0) := x"51"; constant sF99D1A97BFDA9B5076280F23CECAAF884FCBA996 : std_logic_vector(7 downto 0) := x"52"; constant s51302044F211B9E83B0E4160532E89D41D26179F : std_logic_vector(7 downto 0) := x"53"; constant sA0E09E1DFA0715EA5072265E84B3B90BDEF4A330
 : std_logic_vector(7 downto 0) := x"54"; constant s98D7FC4F26467AB3B384D5297B7DAA0066EAB130 : std_logic_vector(7 downto 0) := x"55"; constant s57A7C76B0F0C0E6103B6BDE4922267DFC1C6CAC8 : std_logic_vector(7 downto 0) := x"56"; constant sFAEE7C7664BC579F00801F34E53AA70BD65A7874
 : std_logic_vector(7 downto 0) := x"57"; constant s1E153525FB86CE60222E8A7CBAA485AF861B1D74 : std_logic_vector(7 downto 0) := x"58"; constant s27FC1A1F329912801D6E9215F3007A63A8623499 : std_logic_vector(7 downto 0) := x"59"; constant sE312DD9AD97739BDE32B25BD07E6F495A41E9C6F
 : std_logic_vector(7 downto 0) := x"5A"; constant s97161BEE2D29B3E48064B3B437D9507452C8BE43 : std_logic_vector(7 downto 0) := x"5B";  constant s83F243E9AEA0950EEEE87EEFF9FF2B8AA0412294 : std_logic_vector(7 downto 0) := x"5F";  function sC3DBD2E2D5E3454BB5656AA34F64BFD4C61C3377
 (s6058A04FD298967655739A6C56676FA60DAE306B: in std_logic_vector) return std_logic_vector; end ENDAT_ENCODER_pkg; package body ENDAT_ENCODER_pkg is function sC3DBD2E2D5E3454BB5656AA34F64BFD4C61C3377 (s6058A04FD298967655739A6C56676FA60DAE306B: in std_logic_vector
) return std_logic_vector is variable s7CD850FFC99515521745FADBA902AC96D14969CA: std_logic_vector(s6058A04FD298967655739A6C56676FA60DAE306B'RANGE); alias sE8E6372BF4BD2203497CA7A3D999ACB746D3E75F: std_logic_vector(s6058A04FD298967655739A6C56676FA60DAE306B
'REVERSE_RANGE) is s6058A04FD298967655739A6C56676FA60DAE306B; begin for s020F5125771EEEB6F963720A8BB968FCA977AA41 in sE8E6372BF4BD2203497CA7A3D999ACB746D3E75F'RANGE loop s7CD850FFC99515521745FADBA902AC96D14969CA(s020F5125771EEEB6F963720A8BB968FCA977AA41) := 
sE8E6372BF4BD2203497CA7A3D999ACB746D3E75F(s020F5125771EEEB6F963720A8BB968FCA977AA41); end loop; return s7CD850FFC99515521745FADBA902AC96D14969CA; end;  end ENDAT_ENCODER_pkg; 