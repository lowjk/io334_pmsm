library IEEE; use IEEE.std_logic_1164.all; use IEEE.numeric_std.all; entity PWM_TRIGGER is port ( s82C78E3CD667612DE97ED7C5FA8365F21045093F : in std_logic; s0A61EC3B284D41A7527B973B71395AF396BD0749 : in std_logic; s4F9EF0C7BB9149A40FBFAFB249E3995FB864917A
 : in std_logic; s67BC8086A3CA80A76AC4A164873CAD71C96B5FE0 : in std_logic_vector(7 downto 0); s96088CC8D215E1C4E6BD73028628BBAFD1FB4AB8 : in std_logic_vector(31 downto 0); s160C88F52FE0264EE39CE02AD36940648A499C69 : in std_logic_vector(15 downto 0);  s37394BFF31F8165BDF20DEB888AECA974BBA3623
 : in std_logic_vector(31 downto 0); sBAF99F5E379DD83C7801574B6C9B3543793DAC97 : in std_logic_vector(31 downto 0); s210E8B1235B722AEADE3A804D3F0ABBF1ECDF813 : in std_logic_vector(31 downto 0); s3539C3439A2E15C9F92A30B0F8C66085F38548A7 : in std_logic_vector
(31 downto 0); s176765D58EB0F4B63A08449CD9D42334FA44A80B : in std_logic_vector(31 downto 0); sFEE2B98E596E164B80FA91ED23A3B076B9EF6553 : in std_logic_vector(31 downto 0); sD570C51C1637403B1D115AC1158C653C42ECE9CB : out std_logic ); end PWM_TRIGGER; architecture
 rtl of PWM_TRIGGER is type sA564510C7FCE7940D7D16C6D98FB4EC28EF9532B is (s4CFA0881397DB6939A21DB53B7C9B34BAAD20843, sB8BCC80347362243B5D4480379AC15E39C4DAB51); signal s0FEC712F765FB8844B3F2BBB11D39CEF1DC96CC4, s8E8B32351634161B9B1D8D18043D6DD1583B3BE6 : 
sA564510C7FCE7940D7D16C6D98FB4EC28EF9532B; signal s88E4852E33180732DEC9DF6F65F0A378D208FECF : std_logic; signal s0597C0A28BB30D229FEC515561F1AD824D20604B, sE83A15ECA18BC49D55EB8DDDA31231F41FD522E7 : unsigned(15 downto 0); signal sB8FC36A4D05272CABCCBD52068545D156D0EB94F
 : std_logic; signal s4E1F2C3920D3204BF4351D15F8A4B1EC68E8AF62 : std_logic; begin s88E4852E33180732DEC9DF6F65F0A378D208FECF <= '0' when s4F9EF0C7BB9149A40FBFAFB249E3995FB864917A = '0' else '1' when s67BC8086A3CA80A76AC4A164873CAD71C96B5FE0(0) = '1' and s96088CC8D215E1C4E6BD73028628BBAFD1FB4AB8
 = s37394BFF31F8165BDF20DEB888AECA974BBA3623 else '1' when s67BC8086A3CA80A76AC4A164873CAD71C96B5FE0(1) = '1' and s96088CC8D215E1C4E6BD73028628BBAFD1FB4AB8 = sBAF99F5E379DD83C7801574B6C9B3543793DAC97 else '1' when s67BC8086A3CA80A76AC4A164873CAD71C96B5FE0
(2) = '1' and s96088CC8D215E1C4E6BD73028628BBAFD1FB4AB8 = s210E8B1235B722AEADE3A804D3F0ABBF1ECDF813 else '1' when s67BC8086A3CA80A76AC4A164873CAD71C96B5FE0(3) = '1' and s96088CC8D215E1C4E6BD73028628BBAFD1FB4AB8 = s3539C3439A2E15C9F92A30B0F8C66085F38548A7 
else '1' when s67BC8086A3CA80A76AC4A164873CAD71C96B5FE0(4) = '1' and s96088CC8D215E1C4E6BD73028628BBAFD1FB4AB8 = s176765D58EB0F4B63A08449CD9D42334FA44A80B else '1' when s67BC8086A3CA80A76AC4A164873CAD71C96B5FE0(5) = '1' and s96088CC8D215E1C4E6BD73028628BBAFD1FB4AB8
 = sFEE2B98E596E164B80FA91ED23A3B076B9EF6553 else '0'; process(s0FEC712F765FB8844B3F2BBB11D39CEF1DC96CC4, s88E4852E33180732DEC9DF6F65F0A378D208FECF, s0597C0A28BB30D229FEC515561F1AD824D20604B, s160C88F52FE0264EE39CE02AD36940648A499C69) begin sD570C51C1637403B1D115AC1158C653C42ECE9CB
 <= '0'; sB8FC36A4D05272CABCCBD52068545D156D0EB94F <= '0'; s4E1F2C3920D3204BF4351D15F8A4B1EC68E8AF62 <= '0'; case s0FEC712F765FB8844B3F2BBB11D39CEF1DC96CC4 is when s4CFA0881397DB6939A21DB53B7C9B34BAAD20843 => if s88E4852E33180732DEC9DF6F65F0A378D208FECF = '1' 
then s4E1F2C3920D3204BF4351D15F8A4B1EC68E8AF62 <= '1'; s8E8B32351634161B9B1D8D18043D6DD1583B3BE6 <= sB8BCC80347362243B5D4480379AC15E39C4DAB51; else s8E8B32351634161B9B1D8D18043D6DD1583B3BE6 <= s4CFA0881397DB6939A21DB53B7C9B34BAAD20843; end if; when sB8BCC80347362243B5D4480379AC15E39C4DAB51
 => sD570C51C1637403B1D115AC1158C653C42ECE9CB <= '1'; if s88E4852E33180732DEC9DF6F65F0A378D208FECF = '1' then s4E1F2C3920D3204BF4351D15F8A4B1EC68E8AF62 <= '1'; s8E8B32351634161B9B1D8D18043D6DD1583B3BE6 <= sB8BCC80347362243B5D4480379AC15E39C4DAB51; elsif s0597C0A28BB30D229FEC515561F1AD824D20604B
 = unsigned(s160C88F52FE0264EE39CE02AD36940648A499C69) then s4E1F2C3920D3204BF4351D15F8A4B1EC68E8AF62 <= '1'; s8E8B32351634161B9B1D8D18043D6DD1583B3BE6 <= s4CFA0881397DB6939A21DB53B7C9B34BAAD20843; else sB8FC36A4D05272CABCCBD52068545D156D0EB94F <= '1'; s8E8B32351634161B9B1D8D18043D6DD1583B3BE6
 <= sB8BCC80347362243B5D4480379AC15E39C4DAB51; end if; end case; end process; process(s82C78E3CD667612DE97ED7C5FA8365F21045093F, s0A61EC3B284D41A7527B973B71395AF396BD0749) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749 = '1' then s0FEC712F765FB8844B3F2BBB11D39CEF1DC96CC4
 <= s4CFA0881397DB6939A21DB53B7C9B34BAAD20843; elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then s0FEC712F765FB8844B3F2BBB11D39CEF1DC96CC4 <= s8E8B32351634161B9B1D8D18043D6DD1583B3BE6; end if; end process; process(s82C78E3CD667612DE97ED7C5FA8365F21045093F
, s0A61EC3B284D41A7527B973B71395AF396BD0749) begin if s0A61EC3B284D41A7527B973B71395AF396BD0749 = '1' then s0597C0A28BB30D229FEC515561F1AD824D20604B <= (others => '0'); elsif rising_edge(s82C78E3CD667612DE97ED7C5FA8365F21045093F) then s0597C0A28BB30D229FEC515561F1AD824D20604B
 <= sE83A15ECA18BC49D55EB8DDDA31231F41FD522E7; end if; end process; sE83A15ECA18BC49D55EB8DDDA31231F41FD522E7 <= (others => '0') when s4E1F2C3920D3204BF4351D15F8A4B1EC68E8AF62 = '1' else s0597C0A28BB30D229FEC515561F1AD824D20604B + 1 when sB8FC36A4D05272CABCCBD52068545D156D0EB94F
 = '1' else s0597C0A28BB30D229FEC515561F1AD824D20604B; end rtl;