library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.Numeric_Std.all;
use work.QAE_pkg.all;

entity QAE is
  port(
	  clk_i           : in std_logic; 
    reset_i         : in std_logic; 
    
    version_o       : out std_logic_vector(31 downto 0); 
    
		enable_i        : in std_logic; 
		freeWheel_i     : in std_logic; 
		loadDelta_i     : in std_logic;  
    loadSeg_i       : in std_logic;  
		numSeg_i        : in std_logic_vector(31 downto 0);  
		consign_i       : in std_logic_vector(31 downto 0);  
    delta_i         : in std_logic_vector(31 downto 0);  
    loadDeltaValA_i : in std_logic_vector(31 downto 0);  
    loadDeltaValB_i : in std_logic_vector(31 downto 0);  
    loadSegValA_i   : in std_logic_vector(31 downto 0);  
    loadSegValB_i   : in std_logic_vector(31 downto 0);  
    pos_o           : out std_logic_vector(31 downto 0); 
    a_o             : out std_logic; 
    b_o             : out std_logic; 
    c_o             : out std_logic  
  );
end QAE;

architecture struct of QAE is signal s7BBA3C8AB08CE6CA89340ABD6C98D97CE084FAE3 : std_logic; signal s2C93BAEB1B4BD78658067CD4319B8DDE32E4D483 : std_logic_vector(31 downto 0); begin s6CAE423164E366CDD53B2F8228603558D1938453: entity work.QAE_WHEEL port map( 
s0A61EC3B284D41A7527B973B71395AF396BD0749 => reset_i, s82C78E3CD667612DE97ED7C5FA8365F21045093F => clk_i, s90724AE20811A4A1CF4892AD6C5DE35913A379E1 => s7BBA3C8AB08CE6CA89340ABD6C98D97CE084FAE3, s7414A94932A534C4C1BDB2FEEB2D3AAB8599B128 => numSeg_i, s86FFCF3D164D03DFB129A26F24B615BBF08CCEE0
 => loadDelta_i, s66F6FE61FB267B4B55A1EB5C5A6B5E3162BAD531 => loadSeg_i, s8D38E157D14189FC928FCE48A38AD20C8195C0DF => delta_i, s01C8CEA8B26FE9C07E6D213208100190F11FFC58 => loadDeltaValA_i, s6D1117A4E480A54AA407D7471ABD9B7E03C9B64E => loadSegValA_i, s1BE22644210E653BD6BF626E4CCDC1B4AE2CA9A2
 => s2C93BAEB1B4BD78658067CD4319B8DDE32E4D483, sBE62482AD40DBA872C7029A26677B647B2ACF668 => a_o ); sA8A5B55668CD2040C7ED4C6DD4329D681BA752F4: entity work.QAE_Wheel port map( s0A61EC3B284D41A7527B973B71395AF396BD0749 => reset_i, s82C78E3CD667612DE97ED7C5FA8365F21045093F
 => clk_i, s90724AE20811A4A1CF4892AD6C5DE35913A379E1 => s7BBA3C8AB08CE6CA89340ABD6C98D97CE084FAE3, s7414A94932A534C4C1BDB2FEEB2D3AAB8599B128 => numSeg_i, s86FFCF3D164D03DFB129A26F24B615BBF08CCEE0 => loadDelta_i, s66F6FE61FB267B4B55A1EB5C5A6B5E3162BAD531 => 
loadSeg_i, s8D38E157D14189FC928FCE48A38AD20C8195C0DF => delta_i, s01C8CEA8B26FE9C07E6D213208100190F11FFC58 => loadDeltaValB_i, s6D1117A4E480A54AA407D7471ABD9B7E03C9B64E => loadSegValB_i, s1BE22644210E653BD6BF626E4CCDC1B4AE2CA9A2 => open, sBE62482AD40DBA872C7029A26677B647B2ACF668
 => b_o ); s6586619FAEE639F45226E1515B1E3A4F181407F8: entity work.QAE_POSITIONNER port map( s2BE12327C739923A0BDA5AD372381D3F992B6A0F => s2C93BAEB1B4BD78658067CD4319B8DDE32E4D483, s90724AE20811A4A1CF4892AD6C5DE35913A379E1 => enable_i, s8EC1CD656701F1799C089F63518E2F895FE6470D
 => freeWheel_i, sDF13852084C1BE285B56723469BE3ADFFCF3653B => consign_i, sE3594CA1813735566777C0F293E54987EE6AC901 => s7BBA3C8AB08CE6CA89340ABD6C98D97CE084FAE3 ); version_o <= "10" & s731A256AA7EC109FE962BF102445534C5772925D & s7EC4167F3F7F1E99D074313BF18FF4BA05E7ED10
 & s5907A17D8E29C7EB61D4F347241BFE4DAC407AEA; c_o <= '1' when s2C93BAEB1B4BD78658067CD4319B8DDE32E4D483 = x"00000000" else '0'; pos_o <= s2C93BAEB1B4BD78658067CD4319B8DDE32E4D483; end struct; 